LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
ENTITY TESTBENCH IS
END ENTITY TESTBENCH;
ARCHITECTURE TEST OF TESTBENCH IS
SIGNAL CLOCK_50,RESET,LOAD_CODIFICA,block_sent,UART_TXD,UART_RXD:STD_LOGIC;  
SIGNAL F,T,S,R:STD_LOGIC;
SIGNAL FREQUENZA:STD_LOGIC_VECTOR(3 DOWNTO 0);
SIGNAL PATTERN:STD_LOGIC_VECTOR(7 DOWNTO 0); 
SIGNAL input_codifica:std_logic_vector(15 downto 0); 
  
COMPONENT DUT_HANDLER IS
PORT(
  CLOCK_50,RESET:BUFFER STD_LOGIC;
  load_codifica:buffer std_logic;
  INPUT_CODIFICA: OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
  block_sent,UART_RXD:in std_logic;
  UART_TXD: OUT STD_LOGIC
);  
END COMPONENT; 

COMPONENT pc_interface IS
	PORT 
		(clock, rst_as: IN STD_LOGIC;
		input_codifica: IN STD_LOGIC_VECTOR (15 DOWNTO 0);
		load_codifica: IN STD_LOGIC;
		block_sent: BUFFER STD_LOGIC;
		UART_RXD: IN STD_LOGIC;
		UART_TXD: OUT STD_LOGIC;
		start_ack,read_ack: IN STD_LOGIC;
		F, T, S, R: OUT STD_LOGIC;
		frequenza: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		pattern: OUT STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

BEGIN
  
gestore_dut:DUT_HANDLER port map(CLOCK_50,RESET,LOAD_CODIFICA,INPUT_CODIFICA,block_sent,UART_TXD,UART_RXD);

dut:pc_interface port map
(CLOCK_50,RESET,INPUT_CODIFICA,LOAD_CODIFICA,block_sent,UART_RXD,UART_TXD,'0','0',F,T,S,R,FREQUENZA,PATTERN);  

  
END TEST;