    Mac OS X            	   2  �     �                                    ATTR     �   �   I                  �   9  com.apple.quarantine    �     com.apple.lastuseddate#PS 50-0083;5a5feece;Safari;65639066-4FE9-4750-A56A-50301E6493A9��_Z    ��*#                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          This resource fork intentionally left blank                                                                                                                                                                                                                            ��