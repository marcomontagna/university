XSym
0053
7ba957787278e9540a4df4e0569f9687
/software/dk/nangate45/lef/NangateOpenCellLibrary.lef
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                          