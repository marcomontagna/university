    Mac OS X            	   2  �     �                                    ATTR     �     x                      com.apple.TextEncoding          com.apple.lastuseddate#PS      '   Y  7com.apple.metadata:kMDLabel_4pzwqrpvdq2uidy5xryshnv67u   utf-8;134217984r�`Z    ��<    �roFǹ�~-F`����)�M�k����䍐�Jt��֤��U0�&�|�^�*��:"N�M�� x�����E�A�!h                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                               This resource fork intentionally left blank                                                                                                                                                                                                                            ��