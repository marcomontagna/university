LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
ENTITY TRI_STATE IS
GENERIC (N:INTEGER);
PORT(
ENABLE_OUTPUT	: IN STD_LOGIC;	--segnale di enable, reset e clock
DATA_IN	:	IN STD_LOGIC_VECTOR((N-1) DOWNTO 0);	--dato in ingresso
DATA_OUT	:	OUT STD_LOGIC_VECTOR((N-1) DOWNTO 0) --dato in uscita
);
END ENTITY TRI_STATE;
ARCHITECTURE BEHAVIOR OF TRI_STATE IS
BEGIN
WITH ENABLE_OUTPUT SELECT DATA_OUT<=
DATA_IN WHEN '1',
(OTHERS=>'Z') WHEN OTHERS;
END BEHAVIOR;