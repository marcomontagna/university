LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
ENTITY FLIP_FLOP_D IS
PORT(
EN_REG,CLK,RESET	: IN STD_LOGIC;	--segnale di enable, reset e clock
DATA_REG_IN	:	IN STD_LOGIC;	--dato in ingresso
DATA_REG_OUT	:	OUT STD_LOGIC --dato in uscita
);
END ENTITY FLIP_FLOP_D;
ARCHITECTURE BEHAVIOR OF FLIP_FLOP_D IS
BEGIN
REG_PROCESS: PROCESS(CLK)
BEGIN
IF (CLK'EVENT AND CLK='1') THEN
IF RESET='0' THEN
DATA_REG_OUT<='0';
ELSIF (EN_REG='1') THEN
DATA_REG_OUT<=DATA_REG_IN;
END IF;
END IF;
END PROCESS;
END BEHAVIOR;