
module RCA_GEN_NBIT4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module PGnet_18 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_17 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_16 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_15 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_14 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_13 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_12 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_11 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_10 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_9 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_8 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_7 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_6 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_5 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_4 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_3 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_2 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_1 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_21 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n8), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
endmodule


module PG_20 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n8), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
endmodule


module PG_15 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n8), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
endmodule


module PG_14 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n8), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
endmodule


module PG_9 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n8), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
endmodule


module PG_8 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n8), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
endmodule


module PG_3 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n8), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
endmodule


module PG_2 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n8), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
endmodule


module PG_34 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;
  tri   P;
  tri   G;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_32 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;
  tri   B;
  tri   D;
  tri   G;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_31 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;
  tri   B;
  tri   D;
  tri   G;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_30 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;
  tri   G;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_29 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;
  tri   B;
  tri   D;
  tri   G;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_28 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;
  tri   A;
  tri   C;
  tri   G;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_27 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;
  tri   A;
  tri   C;
  tri   G;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_22 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_19 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_18 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_17 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_16 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_13 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_11 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_10 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_7 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_6 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_5 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_4 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_1 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n8;

  INV_X1 U1 ( .A(n8), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n8) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n14, n15;

  XOR2_X1 U3 ( .A(Ci), .B(n15), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n15) );
  INV_X1 U1 ( .A(n14), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n15), .B2(Ci), .ZN(n14) );
endmodule


module mux21_generic_NBIT4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n16, n17, n18, n19, n20;

  INV_X1 U1 ( .A(SEL), .ZN(n19) );
  INV_X1 U2 ( .A(n18), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n19), .ZN(n18) );
  INV_X1 U4 ( .A(n20), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n19), .ZN(n20) );
  INV_X1 U6 ( .A(n17), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n19), .ZN(n17) );
  INV_X1 U8 ( .A(n16), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n19), .ZN(n16) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module FA_64 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module mux21_generic_NBIT4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n10;

  INV_X1 U1 ( .A(SEL), .ZN(n7) );
  INV_X1 U2 ( .A(n8), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n7), .ZN(n8) );
  INV_X1 U4 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n7), .ZN(n6) );
  INV_X1 U6 ( .A(n9), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n7), .ZN(n9) );
  INV_X1 U8 ( .A(n10), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n7), .ZN(n10) );
endmodule


module mux21_generic_NBIT4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n10;

  INV_X1 U1 ( .A(SEL), .ZN(n7) );
  INV_X1 U2 ( .A(n8), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n7), .ZN(n8) );
  INV_X1 U4 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n7), .ZN(n6) );
  INV_X1 U6 ( .A(n9), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n7), .ZN(n9) );
  INV_X1 U8 ( .A(n10), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n7), .ZN(n10) );
endmodule


module mux21_generic_NBIT4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n10;

  INV_X1 U1 ( .A(SEL), .ZN(n7) );
  INV_X1 U2 ( .A(n8), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n7), .ZN(n8) );
  INV_X1 U4 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n7), .ZN(n6) );
  INV_X1 U6 ( .A(n9), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n7), .ZN(n9) );
  INV_X1 U8 ( .A(n10), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n7), .ZN(n10) );
endmodule


module mux21_generic_NBIT4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n10;

  INV_X1 U1 ( .A(SEL), .ZN(n7) );
  INV_X1 U2 ( .A(n8), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n7), .ZN(n8) );
  INV_X1 U4 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n7), .ZN(n6) );
  INV_X1 U6 ( .A(n9), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n7), .ZN(n9) );
  INV_X1 U8 ( .A(n10), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n7), .ZN(n10) );
endmodule


module mux21_generic_NBIT4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n10;

  INV_X1 U1 ( .A(SEL), .ZN(n7) );
  INV_X1 U2 ( .A(n8), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n7), .ZN(n8) );
  INV_X1 U4 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n7), .ZN(n6) );
  INV_X1 U6 ( .A(n9), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n7), .ZN(n9) );
  INV_X1 U8 ( .A(n10), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n7), .ZN(n10) );
endmodule


module RCA_GEN_NBIT4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21_generic_NBIT4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n7, n8, n9, n10;

  INV_X1 U1 ( .A(SEL), .ZN(n7) );
  INV_X1 U2 ( .A(n8), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n7), .ZN(n8) );
  INV_X1 U4 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U5 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n7), .ZN(n6) );
  INV_X1 U6 ( .A(n9), .ZN(Y[1]) );
  AOI22_X1 U7 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n7), .ZN(n9) );
  INV_X1 U8 ( .A(n10), .ZN(Y[0]) );
  AOI22_X1 U9 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n7), .ZN(n10) );
endmodule


module RCA_GEN_NBIT4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module mux21_generic_NBIT4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;
  wire   n6, n8, n9, n10, n7;

  INV_X1 U1 ( .A(n6), .ZN(Y[3]) );
  AOI22_X1 U2 ( .A1(SEL), .A2(A[3]), .B1(B[3]), .B2(n7), .ZN(n6) );
  INV_X1 U3 ( .A(n8), .ZN(Y[2]) );
  AOI22_X1 U4 ( .A1(A[2]), .A2(SEL), .B1(B[2]), .B2(n7), .ZN(n8) );
  INV_X1 U5 ( .A(n9), .ZN(Y[1]) );
  AOI22_X1 U6 ( .A1(A[1]), .A2(SEL), .B1(B[1]), .B2(n7), .ZN(n9) );
  INV_X1 U7 ( .A(n10), .ZN(Y[0]) );
  AOI22_X1 U8 ( .A1(A[0]), .A2(SEL), .B1(B[0]), .B2(n7), .ZN(n10) );
  INV_X1 U9 ( .A(SEL), .ZN(n7) );
endmodule


module RCA_GEN_NBIT4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_GEN_NBIT4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_64 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module PG_12 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(G) );
  AND2_X1 U2 ( .A1(B), .A2(A), .ZN(P) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
endmodule


module PGnet_19 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_20 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_21 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PG_23 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n2), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
endmodule


module PG_24 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;

  AOI21_X1 U1 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(G) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PGnet_22 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_23 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module PGnet_0 ( A, B, C, P, G );
  input A, B, C;
  output P, G;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(P) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(G) );
endmodule


module carry_select_N4_1 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  wire   sel;
  wire   [3:0] S0;
  wire   [3:0] S1;
  tri   Cin;

  RCA_GEN_NBIT4_2 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_GEN_NBIT4_1 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  mux21_generic_NBIT4_1 MUX1 ( .A(S0), .B(S1), .SEL(sel), .Y(S) );
  INV_X1 U3 ( .A(Cin), .ZN(sel) );
endmodule


module carry_select_N4_2 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  wire   sel;
  wire   [3:0] S0;
  wire   [3:0] S1;
  tri   Cin;

  RCA_GEN_NBIT4_4 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_GEN_NBIT4_3 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  mux21_generic_NBIT4_2 MUX1 ( .A(S0), .B(S1), .SEL(sel), .Y(S) );
  INV_X1 U3 ( .A(Cin), .ZN(sel) );
endmodule


module carry_select_N4_3 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  wire   sel;
  wire   [3:0] S0;
  wire   [3:0] S1;
  tri   Cin;

  RCA_GEN_NBIT4_6 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_GEN_NBIT4_5 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  mux21_generic_NBIT4_3 MUX1 ( .A(S0), .B(S1), .SEL(sel), .Y(S) );
  INV_X1 U3 ( .A(Cin), .ZN(sel) );
endmodule


module carry_select_N4_4 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  wire   sel;
  wire   [3:0] S0;
  wire   [3:0] S1;
  tri   Cin;

  RCA_GEN_NBIT4_8 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_GEN_NBIT4_7 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  mux21_generic_NBIT4_4 MUX1 ( .A(S0), .B(S1), .SEL(sel), .Y(S) );
  INV_X1 U3 ( .A(Cin), .ZN(sel) );
endmodule


module carry_select_N4_5 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  wire   sel;
  wire   [3:0] S0;
  wire   [3:0] S1;
  tri   Cin;

  RCA_GEN_NBIT4_10 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_GEN_NBIT4_9 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  mux21_generic_NBIT4_5 MUX1 ( .A(S0), .B(S1), .SEL(sel), .Y(S) );
  INV_X1 U3 ( .A(Cin), .ZN(sel) );
endmodule


module carry_select_N4_6 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  wire   sel;
  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_GEN_NBIT4_12 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_GEN_NBIT4_11 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  mux21_generic_NBIT4_6 MUX1 ( .A(S0), .B(S1), .SEL(sel), .Y(S) );
  INV_X1 U3 ( .A(Cin), .ZN(sel) );
endmodule


module carry_select_N4_7 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  wire   sel;
  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_GEN_NBIT4_14 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_GEN_NBIT4_13 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  mux21_generic_NBIT4_7 MUX1 ( .A(S0), .B(S1), .SEL(sel), .Y(S) );
  INV_X1 U3 ( .A(Cin), .ZN(sel) );
endmodule


module carry_select_N4_0 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;
  wire   n6;
  wire   [3:0] S0;
  wire   [3:0] S1;

  RCA_GEN_NBIT4_0 RCA1 ( .A(A), .B(B), .Ci(1'b0), .S(S0) );
  RCA_GEN_NBIT4_15 RCA2 ( .A(A), .B(B), .Ci(1'b1), .S(S1) );
  mux21_generic_NBIT4_0 MUX1 ( .A(S0), .B(S1), .SEL(n6), .Y(S) );
  INV_X1 U3 ( .A(Cin), .ZN(n6) );
endmodule


module PG_25 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;
  tri   A;
  tri   C;

  INV_X1 U1 ( .A(n2), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_26 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;

  tri   A;
  tri   B;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_33 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;
  tri   P;
  tri   G;

  AOI21_X1 U1 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
  INV_X1 U2 ( .A(n2), .ZN(G) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_35 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;
  tri   P;
  tri   G;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n2), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
endmodule


module PG_36 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;
  tri   P;
  tri   G;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n2), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
endmodule


module PG_37 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;
  tri   P;
  tri   G;

  INV_X1 U1 ( .A(n2), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_38 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;
  tri   P;
  tri   G;

  INV_X1 U1 ( .A(n2), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_39 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;
  tri   P;
  tri   G;

  INV_X1 U1 ( .A(n2), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_40 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;
  tri   P;
  tri   G;

  INV_X1 U1 ( .A(n2), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module PG_41 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n2), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
endmodule


module PG_42 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n2), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
endmodule


module PG_43 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;

  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(P) );
  INV_X1 U2 ( .A(n2), .ZN(G) );
  AOI21_X1 U3 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
endmodule


module PG_0 ( A, B, C, D, P, G );
  input A, B, C, D;
  output P, G;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(G) );
  AOI21_X1 U2 ( .B1(D), .B2(A), .A(C), .ZN(n2) );
  AND2_X1 U3 ( .A1(B), .A2(A), .ZN(P) );
endmodule


module sparse_tree_carry_gen_4bits_1 ( A, B, c_in, P, G );
  input [3:0] A;
  input [3:0] B;
  input c_in;
  output P, G;
  wire   n3, n4, n5;
  wire   [3:0] P0;
  wire   [3:0] G0;
  wire   [1:0] G1;
  wire   [1:0] P1;

  XOR2_X1 U6 ( .A(B[0]), .B(A[0]), .Z(P0[0]) );
  PGnet_3 pg1_1 ( .A(A[1]), .B(B[1]), .C(1'b0), .P(P0[1]), .G(G0[1]) );
  PGnet_2 pg1_2 ( .A(A[2]), .B(B[2]), .C(1'b0), .P(P0[2]), .G(G0[2]) );
  PGnet_1 pg1_3 ( .A(A[3]), .B(B[3]), .C(1'b0), .P(P0[3]), .G(G0[3]) );
  PG_3 pg2_0 ( .A(P0[1]), .B(P0[0]), .C(G0[1]), .D(G0[0]), .P(P1[0]), .G(G1[0]) );
  PG_2 pg2_1 ( .A(P0[3]), .B(P0[2]), .C(G0[3]), .D(G0[2]), .P(P1[1]), .G(G1[1]) );
  PG_1 pgg ( .A(P1[1]), .B(P1[0]), .C(G1[1]), .D(G1[0]), .P(P), .G(G) );
  AOI21_X1 U2 ( .B1(B[0]), .B2(A[0]), .A(n4), .ZN(n3) );
  INV_X1 U3 ( .A(n5), .ZN(n4) );
  OAI21_X1 U4 ( .B1(A[0]), .B2(B[0]), .A(c_in), .ZN(n5) );
  INV_X1 U5 ( .A(n3), .ZN(G0[0]) );
endmodule


module sparse_tree_carry_gen_4bits_2 ( A, B, c_in, P, G );
  input [3:0] A;
  input [3:0] B;
  input c_in;
  output P, G;
  wire   n3, n4, n5;
  wire   [3:0] P0;
  wire   [3:0] G0;
  wire   [1:0] G1;
  wire   [1:0] P1;

  XOR2_X1 U6 ( .A(B[0]), .B(A[0]), .Z(P0[0]) );
  PGnet_6 pg1_1 ( .A(A[1]), .B(B[1]), .C(1'b0), .P(P0[1]), .G(G0[1]) );
  PGnet_5 pg1_2 ( .A(A[2]), .B(B[2]), .C(1'b0), .P(P0[2]), .G(G0[2]) );
  PGnet_4 pg1_3 ( .A(A[3]), .B(B[3]), .C(1'b0), .P(P0[3]), .G(G0[3]) );
  PG_6 pg2_0 ( .A(P0[1]), .B(P0[0]), .C(G0[1]), .D(G0[0]), .P(P1[0]), .G(G1[0]) );
  PG_5 pg2_1 ( .A(P0[3]), .B(P0[2]), .C(G0[3]), .D(G0[2]), .P(P1[1]), .G(G1[1]) );
  PG_4 pgg ( .A(P1[1]), .B(P1[0]), .C(G1[1]), .D(G1[0]), .P(P), .G(G) );
  INV_X1 U2 ( .A(n3), .ZN(G0[0]) );
  AOI21_X1 U3 ( .B1(B[0]), .B2(A[0]), .A(n4), .ZN(n3) );
  INV_X1 U4 ( .A(n5), .ZN(n4) );
  OAI21_X1 U5 ( .B1(A[0]), .B2(B[0]), .A(c_in), .ZN(n5) );
endmodule


module sparse_tree_carry_gen_4bits_3 ( A, B, c_in, P, G );
  input [3:0] A;
  input [3:0] B;
  input c_in;
  output P, G;
  wire   n3, n4, n5;
  wire   [3:0] P0;
  wire   [3:0] G0;
  wire   [1:0] G1;
  wire   [1:0] P1;

  XOR2_X1 U6 ( .A(B[0]), .B(A[0]), .Z(P0[0]) );
  PGnet_9 pg1_1 ( .A(A[1]), .B(B[1]), .C(1'b0), .P(P0[1]), .G(G0[1]) );
  PGnet_8 pg1_2 ( .A(A[2]), .B(B[2]), .C(1'b0), .P(P0[2]), .G(G0[2]) );
  PGnet_7 pg1_3 ( .A(A[3]), .B(B[3]), .C(1'b0), .P(P0[3]), .G(G0[3]) );
  PG_9 pg2_0 ( .A(P0[1]), .B(P0[0]), .C(G0[1]), .D(G0[0]), .P(P1[0]), .G(G1[0]) );
  PG_8 pg2_1 ( .A(P0[3]), .B(P0[2]), .C(G0[3]), .D(G0[2]), .P(P1[1]), .G(G1[1]) );
  PG_7 pgg ( .A(P1[1]), .B(P1[0]), .C(G1[1]), .D(G1[0]), .P(P), .G(G) );
  AOI21_X1 U2 ( .B1(B[0]), .B2(A[0]), .A(n4), .ZN(n3) );
  INV_X1 U3 ( .A(n5), .ZN(n4) );
  OAI21_X1 U4 ( .B1(A[0]), .B2(B[0]), .A(c_in), .ZN(n5) );
  INV_X1 U5 ( .A(n3), .ZN(G0[0]) );
endmodule


module sparse_tree_carry_gen_4bits_4 ( A, B, c_in, P, G );
  input [3:0] A;
  input [3:0] B;
  input c_in;
  output P, G;
  wire   n3, n4, n5;
  wire   [3:0] P0;
  wire   [3:0] G0;
  wire   [1:0] G1;
  wire   [1:0] P1;

  XOR2_X1 U6 ( .A(B[0]), .B(A[0]), .Z(P0[0]) );
  PGnet_12 pg1_1 ( .A(A[1]), .B(B[1]), .C(1'b0), .P(P0[1]), .G(G0[1]) );
  PGnet_11 pg1_2 ( .A(A[2]), .B(B[2]), .C(1'b0), .P(P0[2]), .G(G0[2]) );
  PGnet_10 pg1_3 ( .A(A[3]), .B(B[3]), .C(1'b0), .P(P0[3]), .G(G0[3]) );
  PG_12 pg2_0 ( .A(P0[1]), .B(P0[0]), .C(G0[1]), .D(G0[0]), .P(P1[0]), .G(
        G1[0]) );
  PG_11 pg2_1 ( .A(P0[3]), .B(P0[2]), .C(G0[3]), .D(G0[2]), .P(P1[1]), .G(
        G1[1]) );
  PG_10 pgg ( .A(P1[1]), .B(P1[0]), .C(G1[1]), .D(G1[0]), .P(P), .G(G) );
  INV_X1 U2 ( .A(n3), .ZN(G0[0]) );
  AOI21_X1 U3 ( .B1(B[0]), .B2(A[0]), .A(n4), .ZN(n3) );
  INV_X1 U4 ( .A(n5), .ZN(n4) );
  OAI21_X1 U5 ( .B1(A[0]), .B2(B[0]), .A(c_in), .ZN(n5) );
endmodule


module sparse_tree_carry_gen_4bits_5 ( A, B, c_in, P, G );
  input [3:0] A;
  input [3:0] B;
  input c_in;
  output P, G;
  wire   n3, n4, n5;
  wire   [3:0] P0;
  wire   [3:0] G0;
  wire   [1:0] G1;
  wire   [1:0] P1;

  XOR2_X1 U6 ( .A(B[0]), .B(A[0]), .Z(P0[0]) );
  PGnet_15 pg1_1 ( .A(A[1]), .B(B[1]), .C(1'b0), .P(P0[1]), .G(G0[1]) );
  PGnet_14 pg1_2 ( .A(A[2]), .B(B[2]), .C(1'b0), .P(P0[2]), .G(G0[2]) );
  PGnet_13 pg1_3 ( .A(A[3]), .B(B[3]), .C(1'b0), .P(P0[3]), .G(G0[3]) );
  PG_15 pg2_0 ( .A(P0[1]), .B(P0[0]), .C(G0[1]), .D(G0[0]), .P(P1[0]), .G(
        G1[0]) );
  PG_14 pg2_1 ( .A(P0[3]), .B(P0[2]), .C(G0[3]), .D(G0[2]), .P(P1[1]), .G(
        G1[1]) );
  PG_13 pgg ( .A(P1[1]), .B(P1[0]), .C(G1[1]), .D(G1[0]), .P(P), .G(G) );
  AOI21_X1 U2 ( .B1(B[0]), .B2(A[0]), .A(n4), .ZN(n3) );
  INV_X1 U3 ( .A(n5), .ZN(n4) );
  OAI21_X1 U4 ( .B1(A[0]), .B2(B[0]), .A(c_in), .ZN(n5) );
  INV_X1 U5 ( .A(n3), .ZN(G0[0]) );
endmodule


module sparse_tree_carry_gen_4bits_6 ( A, B, c_in, P, G );
  input [3:0] A;
  input [3:0] B;
  input c_in;
  output P, G;
  wire   n3, n4, n5;
  wire   [3:0] P0;
  wire   [3:0] G0;
  wire   [1:0] G1;
  wire   [1:0] P1;

  XOR2_X1 U6 ( .A(B[0]), .B(A[0]), .Z(P0[0]) );
  PGnet_18 pg1_1 ( .A(A[1]), .B(B[1]), .C(1'b0), .P(P0[1]), .G(G0[1]) );
  PGnet_17 pg1_2 ( .A(A[2]), .B(B[2]), .C(1'b0), .P(P0[2]), .G(G0[2]) );
  PGnet_16 pg1_3 ( .A(A[3]), .B(B[3]), .C(1'b0), .P(P0[3]), .G(G0[3]) );
  PG_18 pg2_0 ( .A(P0[1]), .B(P0[0]), .C(G0[1]), .D(G0[0]), .P(P1[0]), .G(
        G1[0]) );
  PG_17 pg2_1 ( .A(P0[3]), .B(P0[2]), .C(G0[3]), .D(G0[2]), .P(P1[1]), .G(
        G1[1]) );
  PG_16 pgg ( .A(P1[1]), .B(P1[0]), .C(G1[1]), .D(G1[0]), .P(P), .G(G) );
  INV_X1 U2 ( .A(n3), .ZN(G0[0]) );
  AOI21_X1 U3 ( .B1(B[0]), .B2(A[0]), .A(n4), .ZN(n3) );
  INV_X1 U4 ( .A(n5), .ZN(n4) );
  OAI21_X1 U5 ( .B1(A[0]), .B2(B[0]), .A(c_in), .ZN(n5) );
endmodule


module sparse_tree_carry_gen_4bits_7 ( A, B, c_in, P, G );
  input [3:0] A;
  input [3:0] B;
  input c_in;
  output P, G;
  wire   n3, n4, n5;
  wire   [3:0] P0;
  wire   [3:0] G0;
  wire   [1:0] G1;
  wire   [1:0] P1;

  XOR2_X1 U6 ( .A(B[0]), .B(A[0]), .Z(P0[0]) );
  PGnet_21 pg1_1 ( .A(A[1]), .B(B[1]), .C(1'b0), .P(P0[1]), .G(G0[1]) );
  PGnet_20 pg1_2 ( .A(A[2]), .B(B[2]), .C(1'b0), .P(P0[2]), .G(G0[2]) );
  PGnet_19 pg1_3 ( .A(A[3]), .B(B[3]), .C(1'b0), .P(P0[3]), .G(G0[3]) );
  PG_21 pg2_0 ( .A(P0[1]), .B(P0[0]), .C(G0[1]), .D(G0[0]), .P(P1[0]), .G(
        G1[0]) );
  PG_20 pg2_1 ( .A(P0[3]), .B(P0[2]), .C(G0[3]), .D(G0[2]), .P(P1[1]), .G(
        G1[1]) );
  PG_19 pgg ( .A(P1[1]), .B(P1[0]), .C(G1[1]), .D(G1[0]), .P(P), .G(G) );
  AOI21_X1 U2 ( .B1(B[0]), .B2(A[0]), .A(n4), .ZN(n3) );
  INV_X1 U3 ( .A(n5), .ZN(n4) );
  OAI21_X1 U4 ( .B1(A[0]), .B2(B[0]), .A(c_in), .ZN(n5) );
  INV_X1 U5 ( .A(n3), .ZN(G0[0]) );
endmodule


module sparse_tree_carry_gen_4bits_0 ( A, B, c_in, P, G );
  input [3:0] A;
  input [3:0] B;
  input c_in;
  output P, G;
  wire   n3, n4, n5;
  wire   [3:0] P0;
  wire   [3:0] G0;
  wire   [1:0] G1;
  wire   [1:0] P1;

  XOR2_X1 U6 ( .A(B[0]), .B(A[0]), .Z(P0[0]) );
  PGnet_0 pg1_1 ( .A(A[1]), .B(B[1]), .C(1'b0), .P(P0[1]), .G(G0[1]) );
  PGnet_23 pg1_2 ( .A(A[2]), .B(B[2]), .C(1'b0), .P(P0[2]), .G(G0[2]) );
  PGnet_22 pg1_3 ( .A(A[3]), .B(B[3]), .C(1'b0), .P(P0[3]), .G(G0[3]) );
  PG_24 pg2_0 ( .A(P0[1]), .B(P0[0]), .C(G0[1]), .D(G0[0]), .P(P1[0]), .G(
        G1[0]) );
  PG_23 pg2_1 ( .A(P0[3]), .B(P0[2]), .C(G0[3]), .D(G0[2]), .P(P1[1]), .G(
        G1[1]) );
  PG_22 pgg ( .A(P1[1]), .B(P1[0]), .C(G1[1]), .D(G1[0]), .P(P), .G(G) );
  INV_X1 U2 ( .A(n3), .ZN(G0[0]) );
  INV_X1 U3 ( .A(n5), .ZN(n4) );
  AOI21_X1 U4 ( .B1(B[0]), .B2(A[0]), .A(n4), .ZN(n3) );
  OAI21_X1 U5 ( .B1(A[0]), .B2(B[0]), .A(c_in), .ZN(n5) );
endmodule


module sum_generator_N32_N_carry4 ( A, B, Ci, Sum );
  input [31:0] A;
  input [31:0] B;
  input [8:0] Ci;
  output [31:0] Sum;


  carry_select_N4_0 CBLOCk_0 ( .A(A[3:0]), .B(B[3:0]), .Cin(Ci[0]), .S(
        Sum[3:0]) );
  carry_select_N4_7 CBLOCk_1 ( .A(A[7:4]), .B(B[7:4]), .Cin(Ci[1]), .S(
        Sum[7:4]) );
  carry_select_N4_6 CBLOCk_2 ( .A(A[11:8]), .B(B[11:8]), .Cin(Ci[2]), .S(
        Sum[11:8]) );
  carry_select_N4_5 CBLOCk_3 ( .A(A[15:12]), .B(B[15:12]), .Cin(Ci[3]), .S(
        Sum[15:12]) );
  carry_select_N4_4 CBLOCk_4 ( .A(A[19:16]), .B(B[19:16]), .Cin(Ci[4]), .S(
        Sum[19:16]) );
  carry_select_N4_3 CBLOCk_5 ( .A(A[23:20]), .B(B[23:20]), .Cin(Ci[5]), .S(
        Sum[23:20]) );
  carry_select_N4_2 CBLOCk_6 ( .A(A[27:24]), .B(B[27:24]), .Cin(Ci[6]), .S(
        Sum[27:24]) );
  carry_select_N4_1 CBLOCk_7 ( .A(A[31:28]), .B(B[31:28]), .Cin(Ci[7]), .S(
        Sum[31:28]) );
endmodule


module sparse_tree_carry_gen_N5 ( A, B, C0, Cout );
  input [31:0] A;
  input [31:0] B;
  output [7:0] Cout;
  input C0;
  wire   \G[1][7] , \G[1][5] , \G[1][3] , \G[0][7] , \G[0][6] , \G[0][5] ,
         \G[0][4] , \G[0][3] , \G[0][2] , \G[0][1] , \P[1][7] , \P[1][5] ,
         \P[1][3] , \P[1][1] , \P[1][0] , \P[0][7] , \P[0][6] , \P[0][5] ,
         \P[0][4] , \P[0][3] , \P[0][2] , \P[0][1] , n5, n6;
  tri   \G[2][7] ;
  tri   \G[2][6] ;
  tri   \P[2][7] ;
  tri   \P[2][6] ;
  tri   \P[2][3] ;
  tri   \P[2][2] ;
  assign n5 = C0;

  sparse_tree_carry_gen_4bits_0 pg4_0_0 ( .A(A[3:0]), .B(B[3:0]), .c_in(n6), 
        .P(\P[1][0] ), .G(Cout[0]) );
  sparse_tree_carry_gen_4bits_7 pg4_0_1 ( .A(A[7:4]), .B(B[7:4]), .c_in(n6), 
        .P(\P[0][1] ), .G(\G[0][1] ) );
  sparse_tree_carry_gen_4bits_6 pg4_0_2 ( .A(A[11:8]), .B(B[11:8]), .c_in(n6), 
        .P(\P[0][2] ), .G(\G[0][2] ) );
  sparse_tree_carry_gen_4bits_5 pg4_0_3 ( .A(A[15:12]), .B(B[15:12]), .c_in(n6), .P(\P[0][3] ), .G(\G[0][3] ) );
  sparse_tree_carry_gen_4bits_4 pg4_0_4 ( .A(A[19:16]), .B(B[19:16]), .c_in(n6), .P(\P[0][4] ), .G(\G[0][4] ) );
  sparse_tree_carry_gen_4bits_3 pg4_0_5 ( .A(A[23:20]), .B(B[23:20]), .c_in(n6), .P(\P[0][5] ), .G(\G[0][5] ) );
  sparse_tree_carry_gen_4bits_2 pg4_0_6 ( .A(A[27:24]), .B(B[27:24]), .c_in(n6), .P(\P[0][6] ), .G(\G[0][6] ) );
  sparse_tree_carry_gen_4bits_1 pg4_0_7 ( .A(A[31:28]), .B(B[31:28]), .c_in(n6), .P(\P[0][7] ), .G(\G[0][7] ) );
  PG_0 pg1_1_0 ( .A(\P[0][1] ), .B(\P[1][0] ), .C(\G[0][1] ), .D(Cout[0]), .P(
        \P[1][1] ), .G(Cout[1]) );
  PG_43 pg1_1_1 ( .A(\P[0][3] ), .B(\P[0][2] ), .C(\G[0][3] ), .D(\G[0][2] ), 
        .P(\P[1][3] ), .G(\G[1][3] ) );
  PG_42 pg1_1_2 ( .A(\P[0][5] ), .B(\P[0][4] ), .C(\G[0][5] ), .D(\G[0][4] ), 
        .P(\P[1][5] ), .G(\G[1][5] ) );
  PG_41 pg1_1_3 ( .A(\P[0][7] ), .B(\P[0][6] ), .C(\G[0][7] ), .D(\G[0][6] ), 
        .P(\P[1][7] ), .G(\G[1][7] ) );
  PG_40 gen2_2_0_2_1 ( .A(\P[0][2] ), .B(\P[1][1] ), .C(\G[0][2] ), .D(Cout[1]), .P(\P[2][2] ), .G(Cout[2]) );
  PG_39 gen2_2_0_2_2 ( .A(\P[0][2] ), .B(\P[1][0] ), .C(\G[0][2] ), .D(Cout[0]), .P(\P[2][2] ), .G(Cout[2]) );
  PG_38 gen2_2_0_3_1 ( .A(\P[1][3] ), .B(\P[0][2] ), .C(\G[1][3] ), .D(
        \G[0][2] ), .P(\P[2][3] ), .G(Cout[3]) );
  PG_37 gen2_2_0_3_2 ( .A(\P[1][3] ), .B(\P[1][1] ), .C(\G[1][3] ), .D(Cout[1]), .P(\P[2][3] ), .G(Cout[3]) );
  PG_36 gen2_2_1_6_1 ( .A(\P[0][6] ), .B(\P[1][5] ), .C(\G[0][6] ), .D(
        \G[1][5] ), .P(\P[2][6] ), .G(\G[2][6] ) );
  PG_35 gen2_2_1_6_2 ( .A(\P[0][6] ), .B(\P[0][4] ), .C(\G[0][6] ), .D(
        \G[0][4] ), .P(\P[2][6] ), .G(\G[2][6] ) );
  PG_34 gen2_2_1_7_1 ( .A(\P[1][7] ), .B(\P[0][6] ), .C(\G[1][7] ), .D(
        \G[0][6] ), .P(\P[2][7] ), .G(\G[2][7] ) );
  PG_33 gen2_2_1_7_2 ( .A(\P[1][7] ), .B(\P[1][5] ), .C(\G[1][7] ), .D(
        \G[1][5] ), .P(\P[2][7] ), .G(\G[2][7] ) );
  PG_32 gen2_3_0_4_1 ( .A(\P[0][4] ), .B(\P[2][3] ), .C(\G[0][4] ), .D(Cout[3]), .G(Cout[4]) );
  PG_31 gen2_3_0_4_2 ( .A(\P[0][4] ), .B(\P[2][2] ), .C(\G[0][4] ), .D(Cout[2]), .G(Cout[4]) );
  PG_30 gen2_3_0_5_1 ( .A(\P[1][5] ), .B(\P[0][4] ), .C(\G[1][5] ), .D(
        \G[0][4] ), .G(Cout[5]) );
  PG_29 gen2_3_0_5_2 ( .A(\P[1][5] ), .B(\P[2][3] ), .C(\G[1][5] ), .D(Cout[3]), .G(Cout[5]) );
  PG_28 gen2_3_0_6_1 ( .A(\P[2][6] ), .B(\P[1][5] ), .C(\G[2][6] ), .D(
        \G[1][5] ), .G(Cout[6]) );
  PG_27 gen2_3_0_6_2 ( .A(\P[2][6] ), .B(\P[0][4] ), .C(\G[2][6] ), .D(
        \G[0][4] ), .G(Cout[6]) );
  PG_26 gen2_3_0_7_1 ( .A(\P[2][7] ), .B(\P[2][6] ), .C(\G[2][7] ), .D(
        \G[2][6] ), .G(Cout[7]) );
  PG_25 gen2_3_0_7_2 ( .A(\P[2][7] ), .B(\P[1][5] ), .C(\G[2][7] ), .D(
        \G[1][5] ), .G(Cout[7]) );
  BUF_X1 U1 ( .A(n5), .Z(n6) );
endmodule


module SHIFTER_GENERIC_N32_DW_rbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \MR_int[1][31] , \MR_int[1][30] , \MR_int[1][29] , \MR_int[1][28] ,
         \MR_int[1][27] , \MR_int[1][26] , \MR_int[1][25] , \MR_int[1][24] ,
         \MR_int[1][23] , \MR_int[1][22] , \MR_int[1][21] , \MR_int[1][20] ,
         \MR_int[1][19] , \MR_int[1][18] , \MR_int[1][17] , \MR_int[1][16] ,
         \MR_int[1][15] , \MR_int[1][14] , \MR_int[1][13] , \MR_int[1][12] ,
         \MR_int[1][11] , \MR_int[1][10] , \MR_int[1][9] , \MR_int[1][8] ,
         \MR_int[1][7] , \MR_int[1][6] , \MR_int[1][5] , \MR_int[1][4] ,
         \MR_int[1][3] , \MR_int[1][2] , \MR_int[1][1] , \MR_int[1][0] ,
         \MR_int[2][31] , \MR_int[2][30] , \MR_int[2][29] , \MR_int[2][28] ,
         \MR_int[2][27] , \MR_int[2][26] , \MR_int[2][25] , \MR_int[2][24] ,
         \MR_int[2][23] , \MR_int[2][22] , \MR_int[2][21] , \MR_int[2][20] ,
         \MR_int[2][19] , \MR_int[2][18] , \MR_int[2][17] , \MR_int[2][16] ,
         \MR_int[2][15] , \MR_int[2][14] , \MR_int[2][13] , \MR_int[2][12] ,
         \MR_int[2][11] , \MR_int[2][10] , \MR_int[2][9] , \MR_int[2][8] ,
         \MR_int[2][7] , \MR_int[2][6] , \MR_int[2][5] , \MR_int[2][4] ,
         \MR_int[2][3] , \MR_int[2][2] , \MR_int[2][1] , \MR_int[2][0] ,
         \MR_int[3][31] , \MR_int[3][30] , \MR_int[3][29] , \MR_int[3][28] ,
         \MR_int[3][27] , \MR_int[3][26] , \MR_int[3][25] , \MR_int[3][24] ,
         \MR_int[3][23] , \MR_int[3][22] , \MR_int[3][21] , \MR_int[3][20] ,
         \MR_int[3][19] , \MR_int[3][18] , \MR_int[3][17] , \MR_int[3][16] ,
         \MR_int[3][15] , \MR_int[3][14] , \MR_int[3][13] , \MR_int[3][12] ,
         \MR_int[3][11] , \MR_int[3][10] , \MR_int[3][9] , \MR_int[3][8] ,
         \MR_int[3][7] , \MR_int[3][6] , \MR_int[3][5] , \MR_int[3][4] ,
         \MR_int[3][3] , \MR_int[3][2] , \MR_int[3][1] , \MR_int[3][0] ,
         \MR_int[4][31] , \MR_int[4][30] , \MR_int[4][29] , \MR_int[4][28] ,
         \MR_int[4][27] , \MR_int[4][26] , \MR_int[4][25] , \MR_int[4][24] ,
         \MR_int[4][23] , \MR_int[4][22] , \MR_int[4][21] , \MR_int[4][20] ,
         \MR_int[4][19] , \MR_int[4][18] , \MR_int[4][17] , \MR_int[4][16] ,
         \MR_int[4][15] , \MR_int[4][14] , \MR_int[4][13] , \MR_int[4][12] ,
         \MR_int[4][11] , \MR_int[4][10] , \MR_int[4][9] , \MR_int[4][8] ,
         \MR_int[4][7] , \MR_int[4][6] , \MR_int[4][5] , \MR_int[4][4] ,
         \MR_int[4][3] , \MR_int[4][2] , \MR_int[4][1] , \MR_int[4][0] , n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;

  MUX2_X1 M1_4_31 ( .A(\MR_int[4][31] ), .B(\MR_int[4][15] ), .S(n84), .Z(
        B[31]) );
  MUX2_X1 M1_4_30 ( .A(\MR_int[4][30] ), .B(\MR_int[4][14] ), .S(n84), .Z(
        B[30]) );
  MUX2_X1 M1_4_29 ( .A(\MR_int[4][29] ), .B(\MR_int[4][13] ), .S(n84), .Z(
        B[29]) );
  MUX2_X1 M1_4_28 ( .A(\MR_int[4][28] ), .B(\MR_int[4][12] ), .S(n84), .Z(
        B[28]) );
  MUX2_X1 M1_4_27 ( .A(\MR_int[4][27] ), .B(\MR_int[4][11] ), .S(n84), .Z(
        B[27]) );
  MUX2_X1 M1_4_26 ( .A(\MR_int[4][26] ), .B(\MR_int[4][10] ), .S(n84), .Z(
        B[26]) );
  MUX2_X1 M1_4_25 ( .A(\MR_int[4][25] ), .B(\MR_int[4][9] ), .S(n84), .Z(B[25]) );
  MUX2_X1 M1_4_24 ( .A(\MR_int[4][24] ), .B(\MR_int[4][8] ), .S(n84), .Z(B[24]) );
  MUX2_X1 M1_4_23 ( .A(\MR_int[4][23] ), .B(\MR_int[4][7] ), .S(n84), .Z(B[23]) );
  MUX2_X1 M1_4_22 ( .A(\MR_int[4][22] ), .B(\MR_int[4][6] ), .S(n84), .Z(B[22]) );
  MUX2_X1 M1_4_21 ( .A(\MR_int[4][21] ), .B(\MR_int[4][5] ), .S(n83), .Z(B[21]) );
  MUX2_X1 M1_4_20 ( .A(\MR_int[4][20] ), .B(\MR_int[4][4] ), .S(n83), .Z(B[20]) );
  MUX2_X1 M1_4_19 ( .A(\MR_int[4][19] ), .B(\MR_int[4][3] ), .S(n83), .Z(B[19]) );
  MUX2_X1 M1_4_18 ( .A(\MR_int[4][18] ), .B(\MR_int[4][2] ), .S(n83), .Z(B[18]) );
  MUX2_X1 M1_4_17 ( .A(\MR_int[4][17] ), .B(\MR_int[4][1] ), .S(n83), .Z(B[17]) );
  MUX2_X1 M1_4_16 ( .A(\MR_int[4][16] ), .B(\MR_int[4][0] ), .S(n83), .Z(B[16]) );
  MUX2_X1 M1_4_15 ( .A(\MR_int[4][15] ), .B(\MR_int[4][31] ), .S(n83), .Z(
        B[15]) );
  MUX2_X1 M1_4_14 ( .A(\MR_int[4][14] ), .B(\MR_int[4][30] ), .S(n83), .Z(
        B[14]) );
  MUX2_X1 M1_4_13 ( .A(\MR_int[4][13] ), .B(\MR_int[4][29] ), .S(n83), .Z(
        B[13]) );
  MUX2_X1 M1_4_12 ( .A(\MR_int[4][12] ), .B(\MR_int[4][28] ), .S(n83), .Z(
        B[12]) );
  MUX2_X1 M1_4_11 ( .A(\MR_int[4][11] ), .B(\MR_int[4][27] ), .S(n83), .Z(
        B[11]) );
  MUX2_X1 M1_4_10 ( .A(\MR_int[4][10] ), .B(\MR_int[4][26] ), .S(n82), .Z(
        B[10]) );
  MUX2_X1 M1_4_9 ( .A(\MR_int[4][9] ), .B(\MR_int[4][25] ), .S(n82), .Z(B[9])
         );
  MUX2_X1 M1_4_8 ( .A(\MR_int[4][8] ), .B(\MR_int[4][24] ), .S(n82), .Z(B[8])
         );
  MUX2_X1 M1_4_7 ( .A(\MR_int[4][7] ), .B(\MR_int[4][23] ), .S(n82), .Z(B[7])
         );
  MUX2_X1 M1_4_6 ( .A(\MR_int[4][6] ), .B(\MR_int[4][22] ), .S(n82), .Z(B[6])
         );
  MUX2_X1 M1_4_5 ( .A(\MR_int[4][5] ), .B(\MR_int[4][21] ), .S(n82), .Z(B[5])
         );
  MUX2_X1 M1_4_4 ( .A(\MR_int[4][4] ), .B(\MR_int[4][20] ), .S(n82), .Z(B[4])
         );
  MUX2_X1 M1_4_3 ( .A(\MR_int[4][3] ), .B(\MR_int[4][19] ), .S(n82), .Z(B[3])
         );
  MUX2_X1 M1_4_2 ( .A(\MR_int[4][2] ), .B(\MR_int[4][18] ), .S(n82), .Z(B[2])
         );
  MUX2_X1 M1_4_1 ( .A(\MR_int[4][1] ), .B(\MR_int[4][17] ), .S(n82), .Z(B[1])
         );
  MUX2_X1 M1_4_0 ( .A(\MR_int[4][0] ), .B(\MR_int[4][16] ), .S(n82), .Z(B[0])
         );
  MUX2_X1 M1_3_31_0 ( .A(\MR_int[3][31] ), .B(\MR_int[3][7] ), .S(n81), .Z(
        \MR_int[4][31] ) );
  MUX2_X1 M1_3_30_0 ( .A(\MR_int[3][30] ), .B(\MR_int[3][6] ), .S(n81), .Z(
        \MR_int[4][30] ) );
  MUX2_X1 M1_3_29_0 ( .A(\MR_int[3][29] ), .B(\MR_int[3][5] ), .S(n81), .Z(
        \MR_int[4][29] ) );
  MUX2_X1 M1_3_28_0 ( .A(\MR_int[3][28] ), .B(\MR_int[3][4] ), .S(n81), .Z(
        \MR_int[4][28] ) );
  MUX2_X1 M1_3_27_0 ( .A(\MR_int[3][27] ), .B(\MR_int[3][3] ), .S(n81), .Z(
        \MR_int[4][27] ) );
  MUX2_X1 M1_3_26_0 ( .A(\MR_int[3][26] ), .B(\MR_int[3][2] ), .S(n81), .Z(
        \MR_int[4][26] ) );
  MUX2_X1 M1_3_25_0 ( .A(\MR_int[3][25] ), .B(\MR_int[3][1] ), .S(n81), .Z(
        \MR_int[4][25] ) );
  MUX2_X1 M1_3_24_0 ( .A(\MR_int[3][24] ), .B(\MR_int[3][0] ), .S(n81), .Z(
        \MR_int[4][24] ) );
  MUX2_X1 M1_3_23_0 ( .A(\MR_int[3][23] ), .B(\MR_int[3][31] ), .S(n81), .Z(
        \MR_int[4][23] ) );
  MUX2_X1 M1_3_22_0 ( .A(\MR_int[3][22] ), .B(\MR_int[3][30] ), .S(n81), .Z(
        \MR_int[4][22] ) );
  MUX2_X1 M1_3_21_0 ( .A(\MR_int[3][21] ), .B(\MR_int[3][29] ), .S(n80), .Z(
        \MR_int[4][21] ) );
  MUX2_X1 M1_3_20_0 ( .A(\MR_int[3][20] ), .B(\MR_int[3][28] ), .S(n80), .Z(
        \MR_int[4][20] ) );
  MUX2_X1 M1_3_19_0 ( .A(\MR_int[3][19] ), .B(\MR_int[3][27] ), .S(n80), .Z(
        \MR_int[4][19] ) );
  MUX2_X1 M1_3_18_0 ( .A(\MR_int[3][18] ), .B(\MR_int[3][26] ), .S(n80), .Z(
        \MR_int[4][18] ) );
  MUX2_X1 M1_3_17_0 ( .A(\MR_int[3][17] ), .B(\MR_int[3][25] ), .S(n80), .Z(
        \MR_int[4][17] ) );
  MUX2_X1 M1_3_16_0 ( .A(\MR_int[3][16] ), .B(\MR_int[3][24] ), .S(n80), .Z(
        \MR_int[4][16] ) );
  MUX2_X1 M1_3_15_0 ( .A(\MR_int[3][15] ), .B(\MR_int[3][23] ), .S(n80), .Z(
        \MR_int[4][15] ) );
  MUX2_X1 M1_3_14_0 ( .A(\MR_int[3][14] ), .B(\MR_int[3][22] ), .S(n80), .Z(
        \MR_int[4][14] ) );
  MUX2_X1 M1_3_13_0 ( .A(\MR_int[3][13] ), .B(\MR_int[3][21] ), .S(n80), .Z(
        \MR_int[4][13] ) );
  MUX2_X1 M1_3_12_0 ( .A(\MR_int[3][12] ), .B(\MR_int[3][20] ), .S(n80), .Z(
        \MR_int[4][12] ) );
  MUX2_X1 M1_3_11_0 ( .A(\MR_int[3][11] ), .B(\MR_int[3][19] ), .S(n80), .Z(
        \MR_int[4][11] ) );
  MUX2_X1 M1_3_10_0 ( .A(\MR_int[3][10] ), .B(\MR_int[3][18] ), .S(n79), .Z(
        \MR_int[4][10] ) );
  MUX2_X1 M1_3_9_0 ( .A(\MR_int[3][9] ), .B(\MR_int[3][17] ), .S(n79), .Z(
        \MR_int[4][9] ) );
  MUX2_X1 M1_3_8_0 ( .A(\MR_int[3][8] ), .B(\MR_int[3][16] ), .S(n79), .Z(
        \MR_int[4][8] ) );
  MUX2_X1 M1_3_7 ( .A(\MR_int[3][7] ), .B(\MR_int[3][15] ), .S(n79), .Z(
        \MR_int[4][7] ) );
  MUX2_X1 M1_3_6 ( .A(\MR_int[3][6] ), .B(\MR_int[3][14] ), .S(n79), .Z(
        \MR_int[4][6] ) );
  MUX2_X1 M1_3_5 ( .A(\MR_int[3][5] ), .B(\MR_int[3][13] ), .S(n79), .Z(
        \MR_int[4][5] ) );
  MUX2_X1 M1_3_4 ( .A(\MR_int[3][4] ), .B(\MR_int[3][12] ), .S(n79), .Z(
        \MR_int[4][4] ) );
  MUX2_X1 M1_3_3 ( .A(\MR_int[3][3] ), .B(\MR_int[3][11] ), .S(n79), .Z(
        \MR_int[4][3] ) );
  MUX2_X1 M1_3_2 ( .A(\MR_int[3][2] ), .B(\MR_int[3][10] ), .S(n79), .Z(
        \MR_int[4][2] ) );
  MUX2_X1 M1_3_1 ( .A(\MR_int[3][1] ), .B(\MR_int[3][9] ), .S(n79), .Z(
        \MR_int[4][1] ) );
  MUX2_X1 M1_3_0 ( .A(\MR_int[3][0] ), .B(\MR_int[3][8] ), .S(n79), .Z(
        \MR_int[4][0] ) );
  MUX2_X1 M1_2_31_0 ( .A(\MR_int[2][31] ), .B(\MR_int[2][3] ), .S(n78), .Z(
        \MR_int[3][31] ) );
  MUX2_X1 M1_2_30_0 ( .A(\MR_int[2][30] ), .B(\MR_int[2][2] ), .S(n78), .Z(
        \MR_int[3][30] ) );
  MUX2_X1 M1_2_29_0 ( .A(\MR_int[2][29] ), .B(\MR_int[2][1] ), .S(n78), .Z(
        \MR_int[3][29] ) );
  MUX2_X1 M1_2_28_0 ( .A(\MR_int[2][28] ), .B(\MR_int[2][0] ), .S(n78), .Z(
        \MR_int[3][28] ) );
  MUX2_X1 M1_2_27_0 ( .A(\MR_int[2][27] ), .B(\MR_int[2][31] ), .S(n78), .Z(
        \MR_int[3][27] ) );
  MUX2_X1 M1_2_26_0 ( .A(\MR_int[2][26] ), .B(\MR_int[2][30] ), .S(n78), .Z(
        \MR_int[3][26] ) );
  MUX2_X1 M1_2_25_0 ( .A(\MR_int[2][25] ), .B(\MR_int[2][29] ), .S(n78), .Z(
        \MR_int[3][25] ) );
  MUX2_X1 M1_2_24_0 ( .A(\MR_int[2][24] ), .B(\MR_int[2][28] ), .S(n78), .Z(
        \MR_int[3][24] ) );
  MUX2_X1 M1_2_23_0 ( .A(\MR_int[2][23] ), .B(\MR_int[2][27] ), .S(n78), .Z(
        \MR_int[3][23] ) );
  MUX2_X1 M1_2_22_0 ( .A(\MR_int[2][22] ), .B(\MR_int[2][26] ), .S(n78), .Z(
        \MR_int[3][22] ) );
  MUX2_X1 M1_2_21_0 ( .A(\MR_int[2][21] ), .B(\MR_int[2][25] ), .S(n77), .Z(
        \MR_int[3][21] ) );
  MUX2_X1 M1_2_20_0 ( .A(\MR_int[2][20] ), .B(\MR_int[2][24] ), .S(n77), .Z(
        \MR_int[3][20] ) );
  MUX2_X1 M1_2_19_0 ( .A(\MR_int[2][19] ), .B(\MR_int[2][23] ), .S(n77), .Z(
        \MR_int[3][19] ) );
  MUX2_X1 M1_2_18_0 ( .A(\MR_int[2][18] ), .B(\MR_int[2][22] ), .S(n77), .Z(
        \MR_int[3][18] ) );
  MUX2_X1 M1_2_17_0 ( .A(\MR_int[2][17] ), .B(\MR_int[2][21] ), .S(n77), .Z(
        \MR_int[3][17] ) );
  MUX2_X1 M1_2_16_0 ( .A(\MR_int[2][16] ), .B(\MR_int[2][20] ), .S(n77), .Z(
        \MR_int[3][16] ) );
  MUX2_X1 M1_2_15_0 ( .A(\MR_int[2][15] ), .B(\MR_int[2][19] ), .S(n77), .Z(
        \MR_int[3][15] ) );
  MUX2_X1 M1_2_14_0 ( .A(\MR_int[2][14] ), .B(\MR_int[2][18] ), .S(n77), .Z(
        \MR_int[3][14] ) );
  MUX2_X1 M1_2_13_0 ( .A(\MR_int[2][13] ), .B(\MR_int[2][17] ), .S(n77), .Z(
        \MR_int[3][13] ) );
  MUX2_X1 M1_2_12_0 ( .A(\MR_int[2][12] ), .B(\MR_int[2][16] ), .S(n77), .Z(
        \MR_int[3][12] ) );
  MUX2_X1 M1_2_11_0 ( .A(\MR_int[2][11] ), .B(\MR_int[2][15] ), .S(n77), .Z(
        \MR_int[3][11] ) );
  MUX2_X1 M1_2_10_0 ( .A(\MR_int[2][10] ), .B(\MR_int[2][14] ), .S(n76), .Z(
        \MR_int[3][10] ) );
  MUX2_X1 M1_2_9_0 ( .A(\MR_int[2][9] ), .B(\MR_int[2][13] ), .S(n76), .Z(
        \MR_int[3][9] ) );
  MUX2_X1 M1_2_8_0 ( .A(\MR_int[2][8] ), .B(\MR_int[2][12] ), .S(n76), .Z(
        \MR_int[3][8] ) );
  MUX2_X1 M1_2_7_0 ( .A(\MR_int[2][7] ), .B(\MR_int[2][11] ), .S(n76), .Z(
        \MR_int[3][7] ) );
  MUX2_X1 M1_2_6_0 ( .A(\MR_int[2][6] ), .B(\MR_int[2][10] ), .S(n76), .Z(
        \MR_int[3][6] ) );
  MUX2_X1 M1_2_5_0 ( .A(\MR_int[2][5] ), .B(\MR_int[2][9] ), .S(n76), .Z(
        \MR_int[3][5] ) );
  MUX2_X1 M1_2_4_0 ( .A(\MR_int[2][4] ), .B(\MR_int[2][8] ), .S(n76), .Z(
        \MR_int[3][4] ) );
  MUX2_X1 M1_2_3 ( .A(\MR_int[2][3] ), .B(\MR_int[2][7] ), .S(n76), .Z(
        \MR_int[3][3] ) );
  MUX2_X1 M1_2_2 ( .A(\MR_int[2][2] ), .B(\MR_int[2][6] ), .S(n76), .Z(
        \MR_int[3][2] ) );
  MUX2_X1 M1_2_1 ( .A(\MR_int[2][1] ), .B(\MR_int[2][5] ), .S(n76), .Z(
        \MR_int[3][1] ) );
  MUX2_X1 M1_2_0 ( .A(\MR_int[2][0] ), .B(\MR_int[2][4] ), .S(n76), .Z(
        \MR_int[3][0] ) );
  MUX2_X1 M1_1_31_0 ( .A(\MR_int[1][31] ), .B(\MR_int[1][1] ), .S(n70), .Z(
        \MR_int[2][31] ) );
  MUX2_X1 M1_1_30_0 ( .A(\MR_int[1][30] ), .B(\MR_int[1][0] ), .S(n70), .Z(
        \MR_int[2][30] ) );
  MUX2_X1 M1_1_29_0 ( .A(\MR_int[1][29] ), .B(\MR_int[1][31] ), .S(n70), .Z(
        \MR_int[2][29] ) );
  MUX2_X1 M1_1_28_0 ( .A(\MR_int[1][28] ), .B(\MR_int[1][30] ), .S(n70), .Z(
        \MR_int[2][28] ) );
  MUX2_X1 M1_1_27_0 ( .A(\MR_int[1][27] ), .B(\MR_int[1][29] ), .S(n70), .Z(
        \MR_int[2][27] ) );
  MUX2_X1 M1_1_26_0 ( .A(\MR_int[1][26] ), .B(\MR_int[1][28] ), .S(n70), .Z(
        \MR_int[2][26] ) );
  MUX2_X1 M1_1_25_0 ( .A(\MR_int[1][25] ), .B(\MR_int[1][27] ), .S(n70), .Z(
        \MR_int[2][25] ) );
  MUX2_X1 M1_1_24_0 ( .A(\MR_int[1][24] ), .B(\MR_int[1][26] ), .S(n70), .Z(
        \MR_int[2][24] ) );
  MUX2_X1 M1_1_23_0 ( .A(\MR_int[1][23] ), .B(\MR_int[1][25] ), .S(n70), .Z(
        \MR_int[2][23] ) );
  MUX2_X1 M1_1_22_0 ( .A(\MR_int[1][22] ), .B(\MR_int[1][24] ), .S(n70), .Z(
        \MR_int[2][22] ) );
  MUX2_X1 M1_1_21_0 ( .A(\MR_int[1][21] ), .B(\MR_int[1][23] ), .S(n70), .Z(
        \MR_int[2][21] ) );
  MUX2_X1 M1_1_20_0 ( .A(\MR_int[1][20] ), .B(\MR_int[1][22] ), .S(n71), .Z(
        \MR_int[2][20] ) );
  MUX2_X1 M1_1_19_0 ( .A(\MR_int[1][19] ), .B(\MR_int[1][21] ), .S(n71), .Z(
        \MR_int[2][19] ) );
  MUX2_X1 M1_1_18_0 ( .A(\MR_int[1][18] ), .B(\MR_int[1][20] ), .S(n71), .Z(
        \MR_int[2][18] ) );
  MUX2_X1 M1_1_17_0 ( .A(\MR_int[1][17] ), .B(\MR_int[1][19] ), .S(n71), .Z(
        \MR_int[2][17] ) );
  MUX2_X1 M1_1_16_0 ( .A(\MR_int[1][16] ), .B(\MR_int[1][18] ), .S(n71), .Z(
        \MR_int[2][16] ) );
  MUX2_X1 M1_1_15_0 ( .A(\MR_int[1][15] ), .B(\MR_int[1][17] ), .S(n71), .Z(
        \MR_int[2][15] ) );
  MUX2_X1 M1_1_14_0 ( .A(\MR_int[1][14] ), .B(\MR_int[1][16] ), .S(n71), .Z(
        \MR_int[2][14] ) );
  MUX2_X1 M1_1_13_0 ( .A(\MR_int[1][13] ), .B(\MR_int[1][15] ), .S(n71), .Z(
        \MR_int[2][13] ) );
  MUX2_X1 M1_1_12_0 ( .A(\MR_int[1][12] ), .B(\MR_int[1][14] ), .S(n71), .Z(
        \MR_int[2][12] ) );
  MUX2_X1 M1_1_11_0 ( .A(\MR_int[1][11] ), .B(\MR_int[1][13] ), .S(n71), .Z(
        \MR_int[2][11] ) );
  MUX2_X1 M1_1_10_0 ( .A(\MR_int[1][10] ), .B(\MR_int[1][12] ), .S(n71), .Z(
        \MR_int[2][10] ) );
  MUX2_X1 M1_1_9_0 ( .A(\MR_int[1][9] ), .B(\MR_int[1][11] ), .S(n72), .Z(
        \MR_int[2][9] ) );
  MUX2_X1 M1_1_8_0 ( .A(\MR_int[1][8] ), .B(\MR_int[1][10] ), .S(n72), .Z(
        \MR_int[2][8] ) );
  MUX2_X1 M1_1_7_0 ( .A(\MR_int[1][7] ), .B(\MR_int[1][9] ), .S(n72), .Z(
        \MR_int[2][7] ) );
  MUX2_X1 M1_1_6_0 ( .A(\MR_int[1][6] ), .B(\MR_int[1][8] ), .S(n72), .Z(
        \MR_int[2][6] ) );
  MUX2_X1 M1_1_5_0 ( .A(\MR_int[1][5] ), .B(\MR_int[1][7] ), .S(n72), .Z(
        \MR_int[2][5] ) );
  MUX2_X1 M1_1_4_0 ( .A(\MR_int[1][4] ), .B(\MR_int[1][6] ), .S(n72), .Z(
        \MR_int[2][4] ) );
  MUX2_X1 M1_1_3_0 ( .A(\MR_int[1][3] ), .B(\MR_int[1][5] ), .S(n72), .Z(
        \MR_int[2][3] ) );
  MUX2_X1 M1_1_2_0 ( .A(\MR_int[1][2] ), .B(\MR_int[1][4] ), .S(n72), .Z(
        \MR_int[2][2] ) );
  MUX2_X1 M1_1_1 ( .A(\MR_int[1][1] ), .B(\MR_int[1][3] ), .S(n72), .Z(
        \MR_int[2][1] ) );
  MUX2_X1 M1_1_0 ( .A(\MR_int[1][0] ), .B(\MR_int[1][2] ), .S(n72), .Z(
        \MR_int[2][0] ) );
  MUX2_X1 M1_0_31_0 ( .A(A[31]), .B(A[0]), .S(n75), .Z(\MR_int[1][31] ) );
  MUX2_X1 M1_0_30_0 ( .A(A[30]), .B(A[31]), .S(n75), .Z(\MR_int[1][30] ) );
  MUX2_X1 M1_0_29_0 ( .A(A[29]), .B(A[30]), .S(n75), .Z(\MR_int[1][29] ) );
  MUX2_X1 M1_0_28_0 ( .A(A[28]), .B(A[29]), .S(n75), .Z(\MR_int[1][28] ) );
  MUX2_X1 M1_0_27_0 ( .A(A[27]), .B(A[28]), .S(n75), .Z(\MR_int[1][27] ) );
  MUX2_X1 M1_0_26_0 ( .A(A[26]), .B(A[27]), .S(n75), .Z(\MR_int[1][26] ) );
  MUX2_X1 M1_0_25_0 ( .A(A[25]), .B(A[26]), .S(n75), .Z(\MR_int[1][25] ) );
  MUX2_X1 M1_0_24_0 ( .A(A[24]), .B(A[25]), .S(n75), .Z(\MR_int[1][24] ) );
  MUX2_X1 M1_0_23_0 ( .A(A[23]), .B(A[24]), .S(n75), .Z(\MR_int[1][23] ) );
  MUX2_X1 M1_0_22_0 ( .A(A[22]), .B(A[23]), .S(n75), .Z(\MR_int[1][22] ) );
  MUX2_X1 M1_0_21_0 ( .A(A[21]), .B(A[22]), .S(n74), .Z(\MR_int[1][21] ) );
  MUX2_X1 M1_0_20_0 ( .A(A[20]), .B(A[21]), .S(n74), .Z(\MR_int[1][20] ) );
  MUX2_X1 M1_0_19_0 ( .A(A[19]), .B(A[20]), .S(n74), .Z(\MR_int[1][19] ) );
  MUX2_X1 M1_0_18_0 ( .A(A[18]), .B(A[19]), .S(n74), .Z(\MR_int[1][18] ) );
  MUX2_X1 M1_0_17_0 ( .A(A[17]), .B(A[18]), .S(n74), .Z(\MR_int[1][17] ) );
  MUX2_X1 M1_0_16_0 ( .A(A[16]), .B(A[17]), .S(n74), .Z(\MR_int[1][16] ) );
  MUX2_X1 M1_0_15_0 ( .A(A[15]), .B(A[16]), .S(n74), .Z(\MR_int[1][15] ) );
  MUX2_X1 M1_0_14_0 ( .A(A[14]), .B(A[15]), .S(n74), .Z(\MR_int[1][14] ) );
  MUX2_X1 M1_0_13_0 ( .A(A[13]), .B(A[14]), .S(n74), .Z(\MR_int[1][13] ) );
  MUX2_X1 M1_0_12_0 ( .A(A[12]), .B(A[13]), .S(n74), .Z(\MR_int[1][12] ) );
  MUX2_X1 M1_0_11_0 ( .A(A[11]), .B(A[12]), .S(n74), .Z(\MR_int[1][11] ) );
  MUX2_X1 M1_0_10_0 ( .A(A[10]), .B(A[11]), .S(n73), .Z(\MR_int[1][10] ) );
  MUX2_X1 M1_0_9_0 ( .A(A[9]), .B(A[10]), .S(n73), .Z(\MR_int[1][9] ) );
  MUX2_X1 M1_0_8_0 ( .A(A[8]), .B(A[9]), .S(n73), .Z(\MR_int[1][8] ) );
  MUX2_X1 M1_0_7_0 ( .A(A[7]), .B(A[8]), .S(n73), .Z(\MR_int[1][7] ) );
  MUX2_X1 M1_0_6_0 ( .A(A[6]), .B(A[7]), .S(n73), .Z(\MR_int[1][6] ) );
  MUX2_X1 M1_0_5_0 ( .A(A[5]), .B(A[6]), .S(n73), .Z(\MR_int[1][5] ) );
  MUX2_X1 M1_0_4_0 ( .A(A[4]), .B(A[5]), .S(n73), .Z(\MR_int[1][4] ) );
  MUX2_X1 M1_0_3_0 ( .A(A[3]), .B(A[4]), .S(n73), .Z(\MR_int[1][3] ) );
  MUX2_X1 M1_0_2_0 ( .A(A[2]), .B(A[3]), .S(n73), .Z(\MR_int[1][2] ) );
  MUX2_X1 M1_0_1_0 ( .A(A[1]), .B(A[2]), .S(n73), .Z(\MR_int[1][1] ) );
  MUX2_X1 M1_0_0 ( .A(A[0]), .B(A[1]), .S(n73), .Z(\MR_int[1][0] ) );
  BUF_X1 U2 ( .A(SH[3]), .Z(n79) );
  BUF_X1 U3 ( .A(SH[3]), .Z(n80) );
  BUF_X1 U4 ( .A(SH[4]), .Z(n82) );
  BUF_X1 U5 ( .A(SH[4]), .Z(n83) );
  BUF_X1 U6 ( .A(SH[3]), .Z(n81) );
  BUF_X1 U7 ( .A(SH[4]), .Z(n84) );
  CLKBUF_X1 U8 ( .A(SH[0]), .Z(n73) );
  CLKBUF_X1 U9 ( .A(SH[0]), .Z(n74) );
  CLKBUF_X1 U10 ( .A(SH[2]), .Z(n76) );
  CLKBUF_X1 U11 ( .A(SH[2]), .Z(n77) );
  CLKBUF_X1 U12 ( .A(SH[1]), .Z(n71) );
  CLKBUF_X1 U13 ( .A(SH[1]), .Z(n70) );
  CLKBUF_X1 U14 ( .A(SH[0]), .Z(n75) );
  CLKBUF_X1 U15 ( .A(SH[2]), .Z(n78) );
  CLKBUF_X1 U16 ( .A(SH[1]), .Z(n72) );
endmodule


module SHIFTER_GENERIC_N32_DW_lbsh_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] , n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(n84), .Z(
        B[31]) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(n84), .Z(
        B[30]) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(n84), .Z(
        B[29]) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(n84), .Z(
        B[28]) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(n84), .Z(
        B[27]) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(n84), .Z(
        B[26]) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(n84), .Z(B[25]) );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n84), .Z(B[24]) );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(n84), .Z(B[23]) );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S(n84), .Z(B[22]) );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(n83), .Z(B[21]) );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(n83), .Z(B[20]) );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(n83), .Z(B[19]) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n83), .Z(B[18]) );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(n83), .Z(B[17]) );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(n83), .Z(B[16]) );
  MUX2_X1 M0_4_15 ( .A(\ML_int[4][15] ), .B(\ML_int[4][31] ), .S(n83), .Z(
        B[15]) );
  MUX2_X1 M0_4_14 ( .A(\ML_int[4][14] ), .B(\ML_int[4][30] ), .S(n83), .Z(
        B[14]) );
  MUX2_X1 M0_4_13 ( .A(\ML_int[4][13] ), .B(\ML_int[4][29] ), .S(n83), .Z(
        B[13]) );
  MUX2_X1 M0_4_12 ( .A(\ML_int[4][12] ), .B(\ML_int[4][28] ), .S(n83), .Z(
        B[12]) );
  MUX2_X1 M0_4_11 ( .A(\ML_int[4][11] ), .B(\ML_int[4][27] ), .S(n83), .Z(
        B[11]) );
  MUX2_X1 M0_4_10 ( .A(\ML_int[4][10] ), .B(\ML_int[4][26] ), .S(n82), .Z(
        B[10]) );
  MUX2_X1 M0_4_9 ( .A(\ML_int[4][9] ), .B(\ML_int[4][25] ), .S(n82), .Z(B[9])
         );
  MUX2_X1 M0_4_8 ( .A(\ML_int[4][8] ), .B(\ML_int[4][24] ), .S(n82), .Z(B[8])
         );
  MUX2_X1 M0_4_7 ( .A(\ML_int[4][7] ), .B(\ML_int[4][23] ), .S(n82), .Z(B[7])
         );
  MUX2_X1 M0_4_6 ( .A(\ML_int[4][6] ), .B(\ML_int[4][22] ), .S(n82), .Z(B[6])
         );
  MUX2_X1 M0_4_5 ( .A(\ML_int[4][5] ), .B(\ML_int[4][21] ), .S(n82), .Z(B[5])
         );
  MUX2_X1 M0_4_4 ( .A(\ML_int[4][4] ), .B(\ML_int[4][20] ), .S(n82), .Z(B[4])
         );
  MUX2_X1 M0_4_3 ( .A(\ML_int[4][3] ), .B(\ML_int[4][19] ), .S(n82), .Z(B[3])
         );
  MUX2_X1 M0_4_2 ( .A(\ML_int[4][2] ), .B(\ML_int[4][18] ), .S(n82), .Z(B[2])
         );
  MUX2_X1 M0_4_1 ( .A(\ML_int[4][1] ), .B(\ML_int[4][17] ), .S(n82), .Z(B[1])
         );
  MUX2_X1 M0_4_0 ( .A(\ML_int[4][0] ), .B(\ML_int[4][16] ), .S(n82), .Z(B[0])
         );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n81), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n81), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n81), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n81), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n81), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n81), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n81), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(n81), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n81), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n81), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n80), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n80), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n80), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(n80), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n80), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n80), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n80), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n80), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n80), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n80), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n80), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n79), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n79), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n79), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M0_3_7 ( .A(\ML_int[3][7] ), .B(\ML_int[3][31] ), .S(n79), .Z(
        \ML_int[4][7] ) );
  MUX2_X1 M0_3_6 ( .A(\ML_int[3][6] ), .B(\ML_int[3][30] ), .S(n79), .Z(
        \ML_int[4][6] ) );
  MUX2_X1 M0_3_5 ( .A(\ML_int[3][5] ), .B(\ML_int[3][29] ), .S(n79), .Z(
        \ML_int[4][5] ) );
  MUX2_X1 M0_3_4 ( .A(\ML_int[3][4] ), .B(\ML_int[3][28] ), .S(n79), .Z(
        \ML_int[4][4] ) );
  MUX2_X1 M0_3_3 ( .A(\ML_int[3][3] ), .B(\ML_int[3][27] ), .S(n79), .Z(
        \ML_int[4][3] ) );
  MUX2_X1 M0_3_2 ( .A(\ML_int[3][2] ), .B(\ML_int[3][26] ), .S(n79), .Z(
        \ML_int[4][2] ) );
  MUX2_X1 M0_3_1 ( .A(\ML_int[3][1] ), .B(\ML_int[3][25] ), .S(n79), .Z(
        \ML_int[4][1] ) );
  MUX2_X1 M0_3_0 ( .A(\ML_int[3][0] ), .B(\ML_int[3][24] ), .S(n79), .Z(
        \ML_int[4][0] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(n78), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(n78), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n78), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n78), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(n78), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n78), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n78), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n78), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n78), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n78), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(n76), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n76), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n76), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n76), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(n76), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(n76), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(n76), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n76), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n76), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n76), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n76), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n77), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n77), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n77), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n77), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n77), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n77), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n77), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M0_2_3 ( .A(\ML_int[2][3] ), .B(\ML_int[2][31] ), .S(n77), .Z(
        \ML_int[3][3] ) );
  MUX2_X1 M0_2_2 ( .A(\ML_int[2][2] ), .B(\ML_int[2][30] ), .S(n77), .Z(
        \ML_int[3][2] ) );
  MUX2_X1 M0_2_1 ( .A(\ML_int[2][1] ), .B(\ML_int[2][29] ), .S(n77), .Z(
        \ML_int[3][1] ) );
  MUX2_X1 M0_2_0 ( .A(\ML_int[2][0] ), .B(\ML_int[2][28] ), .S(n77), .Z(
        \ML_int[3][0] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n70), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n70), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n70), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n70), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(n70), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(n70), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(n70), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n70), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n70), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n70), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n70), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n71), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n71), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n71), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n71), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n71), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n71), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n71), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(n71), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n71), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n71), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n71), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n72), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n72), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n72), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n72), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n72), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n72), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n72), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n72), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M0_1_1 ( .A(\ML_int[1][1] ), .B(\ML_int[1][31] ), .S(n72), .Z(
        \ML_int[2][1] ) );
  MUX2_X1 M0_1_0 ( .A(\ML_int[1][0] ), .B(\ML_int[1][30] ), .S(n72), .Z(
        \ML_int[2][0] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(n75), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(n75), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n75), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n75), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n75), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n75), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n75), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n75), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n75), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n75), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(n74), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(n74), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(n74), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(n74), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n74), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(n74), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n74), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n74), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(n74), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(n74), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n74), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n73), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n73), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n73), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n73), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n73), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n73), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n73), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n73), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n73), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n73), .Z(\ML_int[1][1] ) );
  MUX2_X1 M0_0_0 ( .A(A[0]), .B(A[31]), .S(n73), .Z(\ML_int[1][0] ) );
  BUF_X1 U2 ( .A(SH[3]), .Z(n79) );
  BUF_X1 U3 ( .A(SH[3]), .Z(n80) );
  BUF_X1 U4 ( .A(SH[4]), .Z(n82) );
  BUF_X1 U5 ( .A(SH[4]), .Z(n83) );
  BUF_X1 U6 ( .A(SH[3]), .Z(n81) );
  BUF_X1 U7 ( .A(SH[4]), .Z(n84) );
  CLKBUF_X1 U8 ( .A(SH[0]), .Z(n73) );
  CLKBUF_X1 U9 ( .A(SH[0]), .Z(n74) );
  CLKBUF_X1 U10 ( .A(SH[2]), .Z(n77) );
  CLKBUF_X1 U11 ( .A(SH[2]), .Z(n76) );
  CLKBUF_X1 U12 ( .A(SH[1]), .Z(n71) );
  CLKBUF_X1 U13 ( .A(SH[1]), .Z(n70) );
  CLKBUF_X1 U14 ( .A(SH[0]), .Z(n75) );
  CLKBUF_X1 U15 ( .A(SH[2]), .Z(n78) );
  CLKBUF_X1 U16 ( .A(SH[1]), .Z(n72) );
endmodule


module SHIFTER_GENERIC_N32_DW_sra_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[31] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43,
         n45, n47, n48, n49, n50, n51, n52, n54, n56, n57, n58, n59, n60, n61,
         n63, n64, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n95, n96, n98, n99, n100, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n119,
         n122, n125, n126, n129, n130, n131, n132, n133, n136, n139, n140,
         n144, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n166, n167, n168,
         n169, n181, n295, n296, n329, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374;
  assign B[31] = \A[31] ;
  assign \A[31]  = A[31];

  NOR2_X2 U2 ( .A1(n346), .A2(SH[3]), .ZN(n71) );
  NOR2_X2 U3 ( .A1(SH[2]), .A2(SH[3]), .ZN(n73) );
  MUX2_X1 U143 ( .A(\A[31] ), .B(A[30]), .S(n51), .Z(n84) );
  AND2_X1 U4 ( .A1(SH[2]), .A2(n159), .ZN(n10) );
  NOR2_X1 U5 ( .A1(SH[0]), .A2(SH[1]), .ZN(n51) );
  INV_X1 U6 ( .A(n353), .ZN(n349) );
  INV_X1 U7 ( .A(n38), .ZN(n6) );
  NAND2_X1 U8 ( .A1(n71), .A2(n349), .ZN(n38) );
  INV_X1 U9 ( .A(n3), .ZN(n41) );
  OAI21_X1 U10 ( .B1(n351), .B2(n107), .A(n58), .ZN(B[16]) );
  OAI21_X1 U11 ( .B1(n350), .B2(n90), .A(n58), .ZN(B[17]) );
  OAI21_X1 U12 ( .B1(n351), .B2(n59), .A(n58), .ZN(B[18]) );
  OAI21_X1 U13 ( .B1(n350), .B2(n39), .A(n58), .ZN(B[19]) );
  OAI21_X1 U14 ( .B1(n351), .B2(n36), .A(n58), .ZN(B[20]) );
  OAI21_X1 U15 ( .B1(n350), .B2(n33), .A(n58), .ZN(B[21]) );
  OAI21_X1 U16 ( .B1(n350), .B2(n27), .A(n58), .ZN(B[22]) );
  OAI21_X1 U17 ( .B1(n351), .B2(n21), .A(n58), .ZN(B[23]) );
  OAI21_X1 U18 ( .B1(n351), .B2(n14), .A(n58), .ZN(B[24]) );
  OAI21_X1 U19 ( .B1(n350), .B2(n4), .A(n58), .ZN(B[25]) );
  OAI21_X1 U20 ( .B1(n352), .B2(n69), .A(n58), .ZN(B[26]) );
  OAI21_X1 U21 ( .B1(n352), .B2(n68), .A(n58), .ZN(B[27]) );
  OAI21_X1 U22 ( .B1(n352), .B2(n67), .A(n58), .ZN(B[28]) );
  BUF_X1 U23 ( .A(n348), .Z(n353) );
  NAND2_X1 U24 ( .A1(n353), .A2(\A[31] ), .ZN(n58) );
  OAI21_X1 U25 ( .B1(n352), .B2(n66), .A(n58), .ZN(B[29]) );
  OAI21_X1 U26 ( .B1(n352), .B2(n57), .A(n58), .ZN(B[30]) );
  INV_X1 U27 ( .A(n100), .ZN(n74) );
  BUF_X1 U28 ( .A(n347), .Z(n351) );
  BUF_X1 U29 ( .A(n347), .Z(n350) );
  BUF_X1 U30 ( .A(n348), .Z(n352) );
  INV_X1 U31 ( .A(n54), .ZN(n48) );
  INV_X1 U32 ( .A(n56), .ZN(n49) );
  INV_X1 U33 ( .A(n50), .ZN(n43) );
  INV_X1 U34 ( .A(n51), .ZN(n45) );
  NAND2_X1 U35 ( .A1(n73), .A2(n349), .ZN(n3) );
  AOI221_X1 U36 ( .B1(n77), .B2(n71), .C1(n78), .C2(n73), .A(n74), .ZN(n21) );
  AOI221_X1 U37 ( .B1(n75), .B2(n71), .C1(n76), .C2(n73), .A(n74), .ZN(n14) );
  AOI221_X1 U38 ( .B1(n70), .B2(n71), .C1(n72), .C2(n73), .A(n74), .ZN(n4) );
  AOI221_X1 U39 ( .B1(n84), .B2(n71), .C1(n79), .C2(n73), .A(n74), .ZN(n69) );
  AOI221_X1 U40 ( .B1(n18), .B2(n71), .C1(n17), .C2(n73), .A(n162), .ZN(n107)
         );
  INV_X1 U41 ( .A(n163), .ZN(n162) );
  AOI22_X1 U42 ( .A1(n104), .A2(n75), .B1(n83), .B2(n76), .ZN(n163) );
  AOI221_X1 U43 ( .B1(n11), .B2(n71), .C1(n9), .C2(n73), .A(n105), .ZN(n90) );
  INV_X1 U44 ( .A(n106), .ZN(n105) );
  AOI22_X1 U45 ( .A1(n104), .A2(n70), .B1(n83), .B2(n72), .ZN(n106) );
  AOI221_X1 U46 ( .B1(n80), .B2(n71), .C1(n31), .C2(n73), .A(n102), .ZN(n59)
         );
  INV_X1 U47 ( .A(n103), .ZN(n102) );
  AOI22_X1 U48 ( .A1(n104), .A2(n84), .B1(n83), .B2(n79), .ZN(n103) );
  AOI221_X1 U49 ( .B1(n78), .B2(n71), .C1(n25), .C2(n73), .A(n98), .ZN(n39) );
  INV_X1 U50 ( .A(n99), .ZN(n98) );
  AOI21_X1 U51 ( .B1(n83), .B2(n77), .A(n85), .ZN(n99) );
  AOI221_X1 U52 ( .B1(n76), .B2(n71), .C1(n18), .C2(n73), .A(n88), .ZN(n36) );
  INV_X1 U53 ( .A(n89), .ZN(n88) );
  AOI21_X1 U54 ( .B1(n83), .B2(n75), .A(n85), .ZN(n89) );
  AOI221_X1 U55 ( .B1(n72), .B2(n71), .C1(n11), .C2(n73), .A(n86), .ZN(n33) );
  INV_X1 U56 ( .A(n87), .ZN(n86) );
  AOI21_X1 U57 ( .B1(n83), .B2(n70), .A(n85), .ZN(n87) );
  AOI221_X1 U58 ( .B1(n79), .B2(n71), .C1(n80), .C2(n73), .A(n81), .ZN(n27) );
  INV_X1 U59 ( .A(n82), .ZN(n81) );
  AOI21_X1 U60 ( .B1(n83), .B2(n84), .A(n85), .ZN(n82) );
  OAI221_X1 U61 ( .B1(n130), .B2(n3), .C1(n67), .C2(n349), .A(n131), .ZN(B[12]) );
  INV_X1 U62 ( .A(n16), .ZN(n130) );
  AOI222_X1 U63 ( .A1(n6), .A2(n17), .B1(n8), .B2(n18), .C1(n10), .C2(n76), 
        .ZN(n131) );
  OAI221_X1 U64 ( .B1(n26), .B2(n3), .C1(n27), .C2(n349), .A(n28), .ZN(B[6])
         );
  AOI222_X1 U65 ( .A1(n6), .A2(n29), .B1(n8), .B2(n30), .C1(n10), .C2(n31), 
        .ZN(n28) );
  OAI221_X1 U66 ( .B1(n13), .B2(n3), .C1(n14), .C2(n349), .A(n15), .ZN(B[8])
         );
  INV_X1 U67 ( .A(n19), .ZN(n13) );
  AOI222_X1 U68 ( .A1(n6), .A2(n16), .B1(n8), .B2(n17), .C1(n10), .C2(n18), 
        .ZN(n15) );
  OAI221_X1 U69 ( .B1(n35), .B2(n3), .C1(n36), .C2(n349), .A(n37), .ZN(B[4])
         );
  AOI222_X1 U70 ( .A1(n6), .A2(n19), .B1(n8), .B2(n16), .C1(n10), .C2(n17), 
        .ZN(n37) );
  OAI221_X1 U71 ( .B1(n32), .B2(n3), .C1(n33), .C2(n349), .A(n34), .ZN(B[5])
         );
  AOI222_X1 U72 ( .A1(n6), .A2(n12), .B1(n8), .B2(n7), .C1(n10), .C2(n9), .ZN(
        n34) );
  OAI221_X1 U73 ( .B1(n20), .B2(n3), .C1(n21), .C2(n349), .A(n22), .ZN(B[7])
         );
  AOI222_X1 U74 ( .A1(n6), .A2(n23), .B1(n8), .B2(n24), .C1(n10), .C2(n25), 
        .ZN(n22) );
  OAI221_X1 U75 ( .B1(n2), .B2(n3), .C1(n4), .C2(n349), .A(n5), .ZN(B[9]) );
  INV_X1 U76 ( .A(n12), .ZN(n2) );
  AOI222_X1 U77 ( .A1(n6), .A2(n7), .B1(n8), .B2(n9), .C1(n10), .C2(n11), .ZN(
        n5) );
  OAI221_X1 U78 ( .B1(n148), .B2(n3), .C1(n69), .C2(n349), .A(n149), .ZN(B[10]) );
  INV_X1 U79 ( .A(n29), .ZN(n148) );
  AOI222_X1 U80 ( .A1(n6), .A2(n30), .B1(n8), .B2(n31), .C1(n10), .C2(n80), 
        .ZN(n149) );
  OAI221_X1 U81 ( .B1(n132), .B2(n3), .C1(n68), .C2(n349), .A(n133), .ZN(B[11]) );
  INV_X1 U82 ( .A(n23), .ZN(n132) );
  AOI222_X1 U83 ( .A1(n6), .A2(n24), .B1(n8), .B2(n25), .C1(n10), .C2(n78), 
        .ZN(n133) );
  OAI221_X1 U84 ( .B1(n115), .B2(n3), .C1(n66), .C2(n349), .A(n116), .ZN(B[13]) );
  INV_X1 U85 ( .A(n7), .ZN(n115) );
  AOI222_X1 U86 ( .A1(n6), .A2(n9), .B1(n8), .B2(n11), .C1(n10), .C2(n72), 
        .ZN(n116) );
  OAI221_X1 U87 ( .B1(n112), .B2(n3), .C1(n57), .C2(n349), .A(n113), .ZN(B[14]) );
  AOI222_X1 U88 ( .A1(n6), .A2(n31), .B1(n8), .B2(n80), .C1(n10), .C2(n79), 
        .ZN(n113) );
  OAI221_X1 U89 ( .B1(n35), .B2(n38), .C1(n107), .C2(n349), .A(n156), .ZN(B[0]) );
  AOI222_X1 U90 ( .A1(n10), .A2(n16), .B1(n41), .B2(n157), .C1(n8), .C2(n19), 
        .ZN(n156) );
  OAI221_X1 U91 ( .B1(n54), .B2(n354), .C1(n56), .C2(n340), .A(n160), .ZN(n157) );
  OAI221_X1 U92 ( .B1(n32), .B2(n38), .C1(n90), .C2(n349), .A(n91), .ZN(B[1])
         );
  AOI222_X1 U93 ( .A1(n10), .A2(n7), .B1(n41), .B2(n92), .C1(n8), .C2(n12), 
        .ZN(n91) );
  OAI221_X1 U94 ( .B1(n43), .B2(n354), .C1(n45), .C2(n181), .A(n95), .ZN(n92)
         );
  INV_X1 U95 ( .A(A[1]), .ZN(n181) );
  OAI221_X1 U96 ( .B1(n108), .B2(n38), .C1(n109), .C2(n3), .A(n110), .ZN(B[15]) );
  INV_X1 U97 ( .A(n25), .ZN(n108) );
  AOI221_X1 U98 ( .B1(n10), .B2(n77), .C1(n8), .C2(n78), .A(n111), .ZN(n110)
         );
  INV_X1 U99 ( .A(n58), .ZN(n111) );
  AOI21_X1 U100 ( .B1(n77), .B2(n73), .A(n114), .ZN(n68) );
  AOI21_X1 U101 ( .B1(n75), .B2(n73), .A(n114), .ZN(n67) );
  INV_X1 U102 ( .A(n112), .ZN(n30) );
  INV_X1 U103 ( .A(n109), .ZN(n24) );
  BUF_X1 U104 ( .A(SH[4]), .Z(n348) );
  AOI221_X1 U105 ( .B1(n50), .B2(A[7]), .C1(n51), .C2(A[6]), .A(n64), .ZN(n26)
         );
  OAI22_X1 U106 ( .A1(n342), .A2(n54), .B1(n356), .B2(n56), .ZN(n64) );
  OAI21_X1 U107 ( .B1(n346), .B2(n374), .A(n100), .ZN(n114) );
  NOR2_X1 U108 ( .A1(n100), .A2(n346), .ZN(n85) );
  AND2_X1 U109 ( .A1(n159), .A2(n346), .ZN(n8) );
  AND2_X1 U110 ( .A1(SH[3]), .A2(n346), .ZN(n83) );
  AOI21_X1 U111 ( .B1(n70), .B2(n73), .A(n114), .ZN(n66) );
  AOI21_X1 U112 ( .B1(n84), .B2(n73), .A(n114), .ZN(n57) );
  NAND2_X1 U113 ( .A1(\A[31] ), .A2(SH[3]), .ZN(n100) );
  INV_X1 U114 ( .A(n296), .ZN(n295) );
  AND2_X1 U115 ( .A1(SH[3]), .A2(n349), .ZN(n159) );
  BUF_X1 U116 ( .A(SH[4]), .Z(n347) );
  NOR2_X1 U117 ( .A1(n345), .A2(SH[1]), .ZN(n50) );
  OAI221_X1 U118 ( .B1(n43), .B2(n373), .C1(n45), .C2(n371), .A(n166), .ZN(n75) );
  AOI22_X1 U119 ( .A1(A[30]), .A2(n48), .B1(\A[31] ), .B2(n49), .ZN(n166) );
  OAI221_X1 U120 ( .B1(n43), .B2(n367), .C1(n45), .C2(n366), .A(n136), .ZN(n78) );
  AOI22_X1 U121 ( .A1(A[25]), .A2(n48), .B1(A[26]), .B2(n49), .ZN(n136) );
  OAI221_X1 U122 ( .B1(n43), .B2(n368), .C1(n45), .C2(n367), .A(n164), .ZN(n76) );
  AOI22_X1 U123 ( .A1(A[26]), .A2(n48), .B1(A[27]), .B2(n49), .ZN(n164) );
  OAI221_X1 U124 ( .B1(n43), .B2(n369), .C1(n45), .C2(n368), .A(n119), .ZN(n72) );
  AOI22_X1 U125 ( .A1(A[27]), .A2(n48), .B1(A[28]), .B2(n49), .ZN(n119) );
  OAI221_X1 U126 ( .B1(n43), .B2(n370), .C1(n45), .C2(n369), .A(n154), .ZN(n79) );
  AOI22_X1 U127 ( .A1(A[28]), .A2(n48), .B1(n372), .B2(n49), .ZN(n154) );
  OAI221_X1 U128 ( .B1(n43), .B2(n364), .C1(n363), .C2(n45), .A(n168), .ZN(n18) );
  AOI22_X1 U129 ( .A1(A[22]), .A2(n48), .B1(A[23]), .B2(n49), .ZN(n168) );
  OAI221_X1 U130 ( .B1(n43), .B2(n365), .C1(n45), .C2(n364), .A(n122), .ZN(n11) );
  AOI22_X1 U131 ( .A1(A[23]), .A2(n48), .B1(A[24]), .B2(n49), .ZN(n122) );
  OAI221_X1 U132 ( .B1(n43), .B2(n366), .C1(n45), .C2(n365), .A(n150), .ZN(n80) );
  AOI22_X1 U133 ( .A1(A[24]), .A2(n48), .B1(A[25]), .B2(n49), .ZN(n150) );
  OAI221_X1 U134 ( .B1(n43), .B2(n358), .C1(n45), .C2(n344), .A(n161), .ZN(n16) );
  AOI22_X1 U135 ( .A1(n359), .A2(n48), .B1(A[15]), .B2(n49), .ZN(n161) );
  OAI221_X1 U136 ( .B1(n43), .B2(n360), .C1(n45), .C2(n358), .A(n129), .ZN(n7)
         );
  AOI22_X1 U137 ( .A1(A[15]), .A2(n48), .B1(A[16]), .B2(n49), .ZN(n129) );
  OAI221_X1 U138 ( .B1(n43), .B2(n329), .C1(n45), .C2(n361), .A(n125), .ZN(n9)
         );
  AOI22_X1 U139 ( .A1(A[19]), .A2(n48), .B1(A[20]), .B2(n49), .ZN(n125) );
  OAI221_X1 U140 ( .B1(n43), .B2(n371), .C1(n45), .C2(n370), .A(n144), .ZN(n77) );
  AOI22_X1 U141 ( .A1(n372), .A2(n48), .B1(A[30]), .B2(n49), .ZN(n144) );
  OAI221_X1 U142 ( .B1(n363), .B2(n43), .C1(n362), .C2(n45), .A(n139), .ZN(n25) );
  AOI22_X1 U144 ( .A1(A[21]), .A2(n48), .B1(A[22]), .B2(n49), .ZN(n139) );
  OAI221_X1 U145 ( .B1(n362), .B2(n43), .C1(n329), .C2(n45), .A(n151), .ZN(n31) );
  AOI22_X1 U146 ( .A1(A[20]), .A2(n48), .B1(A[21]), .B2(n49), .ZN(n151) );
  OAI221_X1 U147 ( .B1(n43), .B2(n356), .C1(n45), .C2(n342), .A(n158), .ZN(n19) );
  AOI22_X1 U148 ( .A1(A[10]), .A2(n48), .B1(A[11]), .B2(n49), .ZN(n158) );
  OAI221_X1 U149 ( .B1(n43), .B2(n357), .C1(n45), .C2(n356), .A(n93), .ZN(n12)
         );
  AOI22_X1 U150 ( .A1(A[11]), .A2(n48), .B1(A[12]), .B2(n49), .ZN(n93) );
  OAI221_X1 U151 ( .B1(n43), .B2(n343), .C1(n45), .C2(n357), .A(n155), .ZN(n29) );
  AOI22_X1 U152 ( .A1(A[12]), .A2(n48), .B1(A[13]), .B2(n49), .ZN(n155) );
  OAI221_X1 U153 ( .B1(n43), .B2(n344), .C1(n45), .C2(n343), .A(n147), .ZN(n23) );
  AOI22_X1 U154 ( .A1(A[13]), .A2(n48), .B1(n359), .B2(n49), .ZN(n147) );
  NAND2_X1 U155 ( .A1(SH[1]), .A2(n345), .ZN(n54) );
  NAND2_X1 U156 ( .A1(SH[0]), .A2(SH[1]), .ZN(n56) );
  OAI221_X1 U157 ( .B1(n26), .B2(n38), .C1(n59), .C2(n349), .A(n60), .ZN(B[2])
         );
  AOI222_X1 U158 ( .A1(n10), .A2(n30), .B1(n41), .B2(n61), .C1(n8), .C2(n29), 
        .ZN(n60) );
  OAI221_X1 U159 ( .B1(n43), .B2(n340), .C1(n45), .C2(n354), .A(n63), .ZN(n61)
         );
  AOI22_X1 U160 ( .A1(n295), .A2(n48), .B1(A[5]), .B2(n49), .ZN(n63) );
  OAI221_X1 U161 ( .B1(n20), .B2(n38), .C1(n39), .C2(n349), .A(n40), .ZN(B[3])
         );
  AOI222_X1 U162 ( .A1(n10), .A2(n24), .B1(n41), .B2(n42), .C1(n8), .C2(n23), 
        .ZN(n40) );
  OAI221_X1 U163 ( .B1(n43), .B2(n296), .C1(n45), .C2(n340), .A(n47), .ZN(n42)
         );
  AOI22_X1 U164 ( .A1(A[5]), .A2(n48), .B1(A[6]), .B2(n49), .ZN(n47) );
  AOI221_X1 U165 ( .B1(n50), .B2(A[16]), .C1(n51), .C2(A[15]), .A(n140), .ZN(
        n109) );
  OAI22_X1 U166 ( .A1(n361), .A2(n54), .B1(n329), .B2(n56), .ZN(n140) );
  AOI22_X1 U167 ( .A1(A[3]), .A2(n48), .B1(n295), .B2(n49), .ZN(n95) );
  INV_X1 U168 ( .A(n126), .ZN(n70) );
  AOI222_X1 U169 ( .A1(n51), .A2(n372), .B1(n50), .B2(A[30]), .C1(SH[1]), .C2(
        \A[31] ), .ZN(n126) );
  AOI221_X1 U170 ( .B1(n50), .B2(A[15]), .C1(n51), .C2(n359), .A(n152), .ZN(
        n112) );
  INV_X1 U171 ( .A(n153), .ZN(n152) );
  AOI22_X1 U172 ( .A1(A[16]), .A2(n48), .B1(A[17]), .B2(n49), .ZN(n153) );
  OAI221_X1 U173 ( .B1(n54), .B2(n329), .C1(n362), .C2(n56), .A(n167), .ZN(n17) );
  AOI22_X1 U174 ( .A1(A[17]), .A2(n50), .B1(A[16]), .B2(n51), .ZN(n167) );
  AOI221_X1 U175 ( .B1(n50), .B2(A[6]), .C1(n51), .C2(A[5]), .A(n96), .ZN(n32)
         );
  OAI22_X1 U176 ( .A1(n355), .A2(n54), .B1(n342), .B2(n56), .ZN(n96) );
  AOI221_X1 U177 ( .B1(n50), .B2(A[5]), .C1(n51), .C2(n295), .A(n169), .ZN(n35) );
  OAI22_X1 U178 ( .A1(n341), .A2(n54), .B1(n355), .B2(n56), .ZN(n169) );
  AOI221_X1 U179 ( .B1(n50), .B2(A[8]), .C1(n51), .C2(A[7]), .A(n52), .ZN(n20)
         );
  OAI22_X1 U180 ( .A1(n356), .A2(n54), .B1(n357), .B2(n56), .ZN(n52) );
  INV_X1 U181 ( .A(A[18]), .ZN(n329) );
  INV_X1 U182 ( .A(A[7]), .ZN(n355) );
  INV_X1 U183 ( .A(A[4]), .ZN(n296) );
  AND2_X1 U184 ( .A1(SH[2]), .A2(SH[3]), .ZN(n104) );
  INV_X1 U185 ( .A(A[3]), .ZN(n340) );
  INV_X1 U186 ( .A(A[6]), .ZN(n341) );
  INV_X1 U187 ( .A(A[8]), .ZN(n342) );
  INV_X1 U188 ( .A(A[11]), .ZN(n343) );
  INV_X1 U189 ( .A(A[12]), .ZN(n344) );
  AOI22_X1 U190 ( .A1(A[1]), .A2(n50), .B1(A[0]), .B2(n51), .ZN(n160) );
  INV_X1 U191 ( .A(SH[0]), .ZN(n345) );
  INV_X1 U192 ( .A(SH[2]), .ZN(n346) );
  INV_X1 U193 ( .A(A[2]), .ZN(n354) );
  INV_X1 U194 ( .A(A[9]), .ZN(n356) );
  INV_X1 U195 ( .A(A[10]), .ZN(n357) );
  INV_X1 U196 ( .A(A[13]), .ZN(n358) );
  INV_X1 U197 ( .A(n360), .ZN(n359) );
  INV_X1 U198 ( .A(A[14]), .ZN(n360) );
  INV_X1 U199 ( .A(A[17]), .ZN(n361) );
  INV_X1 U200 ( .A(A[19]), .ZN(n362) );
  INV_X1 U201 ( .A(A[20]), .ZN(n363) );
  INV_X1 U202 ( .A(A[21]), .ZN(n364) );
  INV_X1 U203 ( .A(A[22]), .ZN(n365) );
  INV_X1 U204 ( .A(A[23]), .ZN(n366) );
  INV_X1 U205 ( .A(A[24]), .ZN(n367) );
  INV_X1 U206 ( .A(A[25]), .ZN(n368) );
  INV_X1 U207 ( .A(A[26]), .ZN(n369) );
  INV_X1 U208 ( .A(A[27]), .ZN(n370) );
  INV_X1 U209 ( .A(A[28]), .ZN(n371) );
  INV_X1 U210 ( .A(n373), .ZN(n372) );
  INV_X1 U211 ( .A(A[29]), .ZN(n373) );
  INV_X1 U212 ( .A(\A[31] ), .ZN(n374) );
endmodule


module SHIFTER_GENERIC_N32_DW_rash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n46, n48, n51, n52, n53, n58, n59, n60, n61, n62, n63, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n108, n114, n117, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n131, n132, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n150, n152,
         n154, n155, n156, n157, n158, n160, n161, n163, n164, n165, n289,
         n290, n304, n327, n328, n348, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396;

  MUX2_X1 U103 ( .A(n75), .B(n58), .S(SH[2]), .Z(n89) );
  NOR2_X1 U3 ( .A1(n369), .A2(SH[2]), .ZN(n76) );
  INV_X1 U4 ( .A(n3), .ZN(n41) );
  NAND2_X1 U5 ( .A1(n72), .A2(n376), .ZN(n3) );
  INV_X1 U6 ( .A(n373), .ZN(n376) );
  INV_X1 U7 ( .A(n38), .ZN(n6) );
  INV_X1 U8 ( .A(n164), .ZN(n52) );
  NAND2_X1 U9 ( .A1(n73), .A2(n376), .ZN(n38) );
  NOR2_X1 U10 ( .A1(n376), .A2(n124), .ZN(n99) );
  INV_X1 U11 ( .A(n124), .ZN(n72) );
  NOR3_X1 U12 ( .A1(n69), .A2(n370), .A3(n368), .ZN(B[27]) );
  NOR2_X1 U13 ( .A1(n369), .A2(n370), .ZN(n147) );
  NOR2_X1 U14 ( .A1(n370), .A2(n31), .ZN(B[21]) );
  NOR2_X1 U15 ( .A1(n371), .A2(n25), .ZN(B[22]) );
  NOR2_X1 U16 ( .A1(n372), .A2(n19), .ZN(B[23]) );
  NOR2_X1 U17 ( .A1(n371), .A2(n35), .ZN(B[20]) );
  NOR2_X1 U18 ( .A1(n371), .A2(n39), .ZN(B[19]) );
  NOR2_X1 U19 ( .A1(n372), .A2(n4), .ZN(B[25]) );
  NOR2_X1 U20 ( .A1(n372), .A2(n80), .ZN(B[17]) );
  NOR2_X1 U21 ( .A1(n370), .A2(n60), .ZN(B[18]) );
  NOR2_X1 U22 ( .A1(n373), .A2(n95), .ZN(B[16]) );
  NOR2_X1 U23 ( .A1(n372), .A2(n13), .ZN(B[24]) );
  NOR2_X1 U24 ( .A1(n371), .A2(n70), .ZN(B[26]) );
  BUF_X1 U25 ( .A(n375), .Z(n370) );
  INV_X1 U26 ( .A(n12), .ZN(n37) );
  INV_X1 U27 ( .A(n2), .ZN(n33) );
  BUF_X1 U28 ( .A(n374), .Z(n373) );
  AND2_X1 U29 ( .A1(n67), .A2(n41), .ZN(B[29]) );
  AND2_X1 U30 ( .A1(n59), .A2(n41), .ZN(B[30]) );
  AND2_X1 U31 ( .A1(n41), .A2(n58), .ZN(B[31]) );
  BUF_X1 U32 ( .A(n374), .Z(n372) );
  BUF_X1 U33 ( .A(n375), .Z(n371) );
  INV_X1 U34 ( .A(n327), .ZN(n328) );
  INV_X1 U35 ( .A(n289), .ZN(n290) );
  OAI222_X1 U36 ( .A1(n327), .A2(n395), .B1(n163), .B2(n396), .C1(n289), .C2(
        n394), .ZN(n67) );
  NOR2_X2 U37 ( .A1(n367), .A2(n368), .ZN(n73) );
  AOI222_X1 U38 ( .A1(n74), .A2(n73), .B1(n68), .B2(n76), .C1(n17), .C2(n72), 
        .ZN(n35) );
  AOI222_X1 U39 ( .A1(n71), .A2(n73), .B1(n67), .B2(n76), .C1(n11), .C2(n72), 
        .ZN(n31) );
  AOI222_X1 U40 ( .A1(n78), .A2(n73), .B1(n59), .B2(n76), .C1(n79), .C2(n72), 
        .ZN(n25) );
  AOI222_X1 U41 ( .A1(n75), .A2(n73), .B1(n58), .B2(n76), .C1(n77), .C2(n72), 
        .ZN(n19) );
  AOI222_X1 U42 ( .A1(n23), .A2(n72), .B1(n77), .B2(n73), .C1(n89), .C2(n368), 
        .ZN(n39) );
  INV_X1 U43 ( .A(n44), .ZN(n51) );
  AOI221_X1 U44 ( .B1(n51), .B2(A[11]), .C1(n52), .C2(A[10]), .A(n146), .ZN(
        n12) );
  OAI22_X1 U45 ( .A1(n379), .A2(n327), .B1(n363), .B2(n289), .ZN(n146) );
  AOI221_X1 U46 ( .B1(n51), .B2(A[12]), .C1(n52), .C2(A[11]), .A(n83), .ZN(n2)
         );
  OAI22_X1 U47 ( .A1(n380), .A2(n327), .B1(n379), .B2(n289), .ZN(n83) );
  AOI221_X1 U48 ( .B1(n17), .B2(n73), .C1(n16), .C2(n72), .A(n154), .ZN(n95)
         );
  INV_X1 U49 ( .A(n155), .ZN(n154) );
  AOI22_X1 U50 ( .A1(n92), .A2(n68), .B1(n76), .B2(n74), .ZN(n155) );
  AOI221_X1 U51 ( .B1(n11), .B2(n73), .C1(n9), .C2(n72), .A(n93), .ZN(n80) );
  INV_X1 U52 ( .A(n94), .ZN(n93) );
  AOI22_X1 U53 ( .A1(n92), .A2(n67), .B1(n76), .B2(n71), .ZN(n94) );
  OAI221_X1 U54 ( .B1(n97), .B2(n38), .C1(n43), .C2(n3), .A(n125), .ZN(B[11])
         );
  AOI221_X1 U55 ( .B1(n10), .B2(n77), .C1(n8), .C2(n23), .A(n126), .ZN(n125)
         );
  NOR3_X1 U56 ( .A1(n376), .A2(n368), .A3(n69), .ZN(n126) );
  INV_X1 U57 ( .A(n121), .ZN(B[12]) );
  AOI221_X1 U58 ( .B1(n16), .B2(n6), .C1(n15), .C2(n41), .A(n122), .ZN(n121)
         );
  INV_X1 U59 ( .A(n123), .ZN(n122) );
  AOI222_X1 U60 ( .A1(n10), .A2(n74), .B1(n99), .B2(n68), .C1(n8), .C2(n17), 
        .ZN(n123) );
  AND2_X1 U61 ( .A1(n147), .A2(n367), .ZN(n8) );
  OAI221_X1 U62 ( .B1(n34), .B2(n3), .C1(n35), .C2(n376), .A(n36), .ZN(B[4])
         );
  AOI222_X1 U63 ( .A1(n6), .A2(n37), .B1(n8), .B2(n15), .C1(n10), .C2(n16), 
        .ZN(n36) );
  OAI221_X1 U64 ( .B1(n30), .B2(n3), .C1(n31), .C2(n376), .A(n32), .ZN(B[5])
         );
  AOI222_X1 U65 ( .A1(n6), .A2(n33), .B1(n8), .B2(n7), .C1(n10), .C2(n9), .ZN(
        n32) );
  OAI221_X1 U66 ( .B1(n24), .B2(n3), .C1(n25), .C2(n376), .A(n26), .ZN(B[6])
         );
  AOI222_X1 U67 ( .A1(n6), .A2(n27), .B1(n8), .B2(n28), .C1(n10), .C2(n29), 
        .ZN(n26) );
  OAI221_X1 U68 ( .B1(n18), .B2(n3), .C1(n19), .C2(n376), .A(n20), .ZN(B[7])
         );
  AOI222_X1 U69 ( .A1(n6), .A2(n21), .B1(n8), .B2(n22), .C1(n10), .C2(n23), 
        .ZN(n20) );
  OAI221_X1 U70 ( .B1(n12), .B2(n3), .C1(n13), .C2(n376), .A(n14), .ZN(B[8])
         );
  AOI222_X1 U71 ( .A1(n6), .A2(n15), .B1(n8), .B2(n16), .C1(n10), .C2(n17), 
        .ZN(n14) );
  OAI221_X1 U72 ( .B1(n2), .B2(n3), .C1(n4), .C2(n376), .A(n5), .ZN(B[9]) );
  AOI222_X1 U73 ( .A1(n6), .A2(n7), .B1(n8), .B2(n9), .C1(n10), .C2(n11), .ZN(
        n5) );
  OAI221_X1 U74 ( .B1(n63), .B2(n3), .C1(n70), .C2(n376), .A(n138), .ZN(B[10])
         );
  AOI222_X1 U75 ( .A1(n6), .A2(n28), .B1(n8), .B2(n29), .C1(n10), .C2(n79), 
        .ZN(n138) );
  OAI221_X1 U76 ( .B1(n34), .B2(n38), .C1(n95), .C2(n376), .A(n144), .ZN(B[0])
         );
  AOI222_X1 U77 ( .A1(n10), .A2(n15), .B1(n41), .B2(n145), .C1(n8), .C2(n37), 
        .ZN(n144) );
  OAI221_X1 U78 ( .B1(n44), .B2(n359), .C1(n163), .C2(n377), .A(n150), .ZN(
        n145) );
  OAI221_X1 U79 ( .B1(n30), .B2(n38), .C1(n80), .C2(n376), .A(n81), .ZN(B[1])
         );
  AOI222_X1 U80 ( .A1(n10), .A2(n7), .B1(n41), .B2(n82), .C1(n8), .C2(n33), 
        .ZN(n81) );
  OAI221_X1 U81 ( .B1(n44), .B2(n304), .C1(n165), .C2(n359), .A(n87), .ZN(n82)
         );
  AOI22_X1 U82 ( .A1(A[2]), .A2(n328), .B1(A[1]), .B2(n290), .ZN(n87) );
  OAI221_X1 U83 ( .B1(n103), .B2(n38), .C1(n104), .C2(n3), .A(n105), .ZN(B[13]) );
  INV_X1 U84 ( .A(n7), .ZN(n104) );
  INV_X1 U85 ( .A(n9), .ZN(n103) );
  AOI222_X1 U86 ( .A1(n10), .A2(n71), .B1(n99), .B2(n67), .C1(n8), .C2(n11), 
        .ZN(n105) );
  OAI221_X1 U87 ( .B1(n100), .B2(n38), .C1(n101), .C2(n3), .A(n102), .ZN(B[14]) );
  INV_X1 U88 ( .A(n28), .ZN(n101) );
  INV_X1 U89 ( .A(n29), .ZN(n100) );
  AOI222_X1 U90 ( .A1(n10), .A2(n78), .B1(n99), .B2(n59), .C1(n8), .C2(n79), 
        .ZN(n102) );
  OAI221_X1 U91 ( .B1(n96), .B2(n38), .C1(n97), .C2(n3), .A(n98), .ZN(B[15])
         );
  INV_X1 U92 ( .A(n23), .ZN(n96) );
  AOI222_X1 U93 ( .A1(n10), .A2(n75), .B1(n99), .B2(n58), .C1(n8), .C2(n77), 
        .ZN(n98) );
  NOR2_X1 U94 ( .A1(n396), .A2(n289), .ZN(n58) );
  AOI22_X1 U95 ( .A1(n74), .A2(n72), .B1(n68), .B2(n73), .ZN(n13) );
  AOI22_X1 U96 ( .A1(n71), .A2(n72), .B1(n67), .B2(n73), .ZN(n4) );
  AOI22_X1 U97 ( .A1(n78), .A2(n72), .B1(n59), .B2(n73), .ZN(n70) );
  BUF_X1 U98 ( .A(n46), .Z(n163) );
  BUF_X1 U99 ( .A(n46), .Z(n164) );
  AOI221_X1 U100 ( .B1(n79), .B2(n73), .C1(n29), .C2(n72), .A(n90), .ZN(n60)
         );
  INV_X1 U101 ( .A(n91), .ZN(n90) );
  AOI22_X1 U102 ( .A1(n92), .A2(n59), .B1(n76), .B2(n78), .ZN(n91) );
  INV_X1 U104 ( .A(SH[3]), .ZN(n369) );
  NAND2_X1 U105 ( .A1(n367), .A2(n369), .ZN(n124) );
  INV_X1 U106 ( .A(n22), .ZN(n97) );
  INV_X1 U107 ( .A(n63), .ZN(n27) );
  INV_X1 U108 ( .A(n43), .ZN(n21) );
  INV_X1 U109 ( .A(n89), .ZN(n69) );
  AND2_X1 U110 ( .A1(n68), .A2(n41), .ZN(B[28]) );
  BUF_X1 U111 ( .A(SH[4]), .Z(n374) );
  BUF_X1 U112 ( .A(SH[4]), .Z(n375) );
  OAI22_X1 U113 ( .A1(n289), .A2(n395), .B1(n327), .B2(n396), .ZN(n59) );
  AOI221_X1 U114 ( .B1(n51), .B2(n362), .C1(n52), .C2(A[7]), .A(n88), .ZN(n30)
         );
  OAI22_X1 U115 ( .A1(n361), .A2(n327), .B1(n360), .B2(n289), .ZN(n88) );
  AOI221_X1 U116 ( .B1(n51), .B2(A[9]), .C1(n52), .C2(n362), .A(n66), .ZN(n24)
         );
  OAI22_X1 U117 ( .A1(n378), .A2(n327), .B1(n361), .B2(n289), .ZN(n66) );
  AOI221_X1 U118 ( .B1(n51), .B2(A[10]), .C1(n52), .C2(A[9]), .A(n53), .ZN(n18) );
  OAI22_X1 U119 ( .A1(n363), .A2(n327), .B1(n378), .B2(n289), .ZN(n53) );
  NOR2_X1 U120 ( .A1(n367), .A2(n369), .ZN(n92) );
  BUF_X1 U121 ( .A(n46), .Z(n165) );
  NAND2_X1 U122 ( .A1(SH[1]), .A2(SH[0]), .ZN(n44) );
  AND2_X1 U123 ( .A1(SH[2]), .A2(n147), .ZN(n10) );
  OR2_X1 U124 ( .A1(SH[0]), .A2(SH[1]), .ZN(n289) );
  OR2_X1 U125 ( .A1(n366), .A2(SH[1]), .ZN(n327) );
  OAI221_X1 U126 ( .B1(n44), .B2(n385), .C1(n164), .C2(n348), .A(n158), .ZN(
        n16) );
  AOI22_X1 U127 ( .A1(A[17]), .A2(n328), .B1(A[16]), .B2(n290), .ZN(n158) );
  OAI221_X1 U128 ( .B1(n44), .B2(n383), .C1(n163), .C2(n382), .A(n117), .ZN(n7) );
  AOI22_X1 U129 ( .A1(A[14]), .A2(n328), .B1(A[13]), .B2(n290), .ZN(n117) );
  OAI221_X1 U130 ( .B1(n44), .B2(n384), .C1(n165), .C2(n383), .A(n141), .ZN(
        n28) );
  AOI22_X1 U131 ( .A1(A[15]), .A2(n328), .B1(A[14]), .B2(n290), .ZN(n141) );
  OAI221_X1 U132 ( .B1(n44), .B2(n382), .C1(n163), .C2(n381), .A(n152), .ZN(
        n15) );
  AOI22_X1 U133 ( .A1(A[13]), .A2(n328), .B1(A[12]), .B2(n290), .ZN(n152) );
  OAI221_X1 U134 ( .B1(n44), .B2(n392), .C1(n164), .C2(n391), .A(n156), .ZN(
        n74) );
  AOI22_X1 U135 ( .A1(A[25]), .A2(n328), .B1(A[24]), .B2(n290), .ZN(n156) );
  OAI221_X1 U136 ( .B1(n44), .B2(n393), .C1(n163), .C2(n392), .A(n114), .ZN(
        n71) );
  AOI22_X1 U137 ( .A1(A[26]), .A2(n328), .B1(A[25]), .B2(n290), .ZN(n114) );
  OAI221_X1 U138 ( .B1(n44), .B2(n389), .C1(n163), .C2(n388), .A(n108), .ZN(
        n11) );
  AOI22_X1 U139 ( .A1(A[22]), .A2(n328), .B1(A[21]), .B2(n290), .ZN(n108) );
  OAI221_X1 U140 ( .B1(n44), .B2(n391), .C1(n164), .C2(n390), .A(n131), .ZN(
        n77) );
  AOI22_X1 U141 ( .A1(A[24]), .A2(n328), .B1(A[23]), .B2(n290), .ZN(n131) );
  OAI221_X1 U142 ( .B1(n386), .B2(n327), .C1(n385), .C2(n289), .A(n128), .ZN(
        n23) );
  AOI22_X1 U143 ( .A1(A[22]), .A2(n51), .B1(A[21]), .B2(n52), .ZN(n128) );
  OAI221_X1 U144 ( .B1(n385), .B2(n327), .C1(n348), .C2(n289), .A(n140), .ZN(
        n29) );
  AOI22_X1 U145 ( .A1(A[21]), .A2(n51), .B1(n52), .B2(A[20]), .ZN(n140) );
  OAI221_X1 U146 ( .B1(n327), .B2(n387), .C1(n386), .C2(n289), .A(n160), .ZN(
        n17) );
  AOI22_X1 U147 ( .A1(A[23]), .A2(n51), .B1(A[22]), .B2(n52), .ZN(n160) );
  OAI221_X1 U148 ( .B1(n44), .B2(n348), .C1(n165), .C2(n384), .A(n137), .ZN(
        n22) );
  AOI22_X1 U149 ( .A1(A[16]), .A2(n328), .B1(A[15]), .B2(n290), .ZN(n137) );
  AOI221_X1 U150 ( .B1(n51), .B2(A[13]), .C1(n52), .C2(A[12]), .A(n143), .ZN(
        n63) );
  OAI22_X1 U151 ( .A1(n364), .A2(n327), .B1(n380), .B2(n289), .ZN(n143) );
  AOI221_X1 U152 ( .B1(n51), .B2(A[14]), .C1(n52), .C2(A[13]), .A(n132), .ZN(
        n43) );
  OAI22_X1 U153 ( .A1(n365), .A2(n327), .B1(n364), .B2(n289), .ZN(n132) );
  OAI221_X1 U154 ( .B1(n44), .B2(n395), .C1(n164), .C2(n394), .A(n127), .ZN(
        n75) );
  AOI22_X1 U155 ( .A1(A[28]), .A2(n328), .B1(A[27]), .B2(n290), .ZN(n127) );
  OAI221_X1 U156 ( .B1(n24), .B2(n38), .C1(n60), .C2(n376), .A(n61), .ZN(B[2])
         );
  AOI222_X1 U157 ( .A1(n10), .A2(n28), .B1(n41), .B2(n62), .C1(n8), .C2(n27), 
        .ZN(n61) );
  OAI221_X1 U158 ( .B1(n44), .B2(n360), .C1(n165), .C2(n304), .A(n65), .ZN(n62) );
  AOI22_X1 U159 ( .A1(A[3]), .A2(n328), .B1(A[2]), .B2(n290), .ZN(n65) );
  OAI221_X1 U160 ( .B1(n18), .B2(n38), .C1(n39), .C2(n376), .A(n40), .ZN(B[3])
         );
  AOI222_X1 U161 ( .A1(n10), .A2(n22), .B1(n41), .B2(n42), .C1(n8), .C2(n21), 
        .ZN(n40) );
  OAI221_X1 U162 ( .B1(n44), .B2(n361), .C1(n165), .C2(n360), .A(n48), .ZN(n42) );
  AOI22_X1 U163 ( .A1(A[4]), .A2(n328), .B1(A[3]), .B2(n290), .ZN(n48) );
  OAI221_X1 U164 ( .B1(n44), .B2(n386), .C1(n164), .C2(n385), .A(n120), .ZN(n9) );
  AOI22_X1 U165 ( .A1(A[18]), .A2(n328), .B1(A[17]), .B2(n290), .ZN(n120) );
  OAI221_X1 U166 ( .B1(n44), .B2(n390), .C1(n165), .C2(n389), .A(n139), .ZN(
        n79) );
  AOI22_X1 U167 ( .A1(A[23]), .A2(n328), .B1(A[22]), .B2(n290), .ZN(n139) );
  OAI221_X1 U168 ( .B1(n44), .B2(n396), .C1(n164), .C2(n395), .A(n157), .ZN(
        n68) );
  AOI22_X1 U169 ( .A1(A[29]), .A2(n328), .B1(A[28]), .B2(n290), .ZN(n157) );
  OAI221_X1 U170 ( .B1(n44), .B2(n394), .C1(n163), .C2(n393), .A(n142), .ZN(
        n78) );
  AOI22_X1 U171 ( .A1(A[27]), .A2(n328), .B1(A[26]), .B2(n290), .ZN(n142) );
  NAND2_X1 U172 ( .A1(SH[1]), .A2(n366), .ZN(n46) );
  AOI221_X1 U173 ( .B1(n51), .B2(A[7]), .C1(n52), .C2(A[6]), .A(n161), .ZN(n34) );
  OAI22_X1 U174 ( .A1(n360), .A2(n327), .B1(n304), .B2(n289), .ZN(n161) );
  INV_X1 U175 ( .A(A[8]), .ZN(n363) );
  INV_X1 U176 ( .A(A[4]), .ZN(n304) );
  INV_X1 U177 ( .A(A[11]), .ZN(n364) );
  INV_X1 U178 ( .A(A[7]), .ZN(n378) );
  INV_X1 U179 ( .A(A[9]), .ZN(n379) );
  INV_X1 U180 ( .A(A[10]), .ZN(n380) );
  INV_X1 U181 ( .A(A[18]), .ZN(n348) );
  INV_X1 U182 ( .A(A[3]), .ZN(n359) );
  INV_X1 U183 ( .A(A[5]), .ZN(n360) );
  INV_X1 U184 ( .A(A[6]), .ZN(n361) );
  INV_X1 U185 ( .A(n363), .ZN(n362) );
  INV_X1 U186 ( .A(A[12]), .ZN(n365) );
  AOI22_X1 U187 ( .A1(A[1]), .A2(n328), .B1(A[0]), .B2(n290), .ZN(n150) );
  INV_X1 U188 ( .A(SH[0]), .ZN(n366) );
  INV_X1 U189 ( .A(SH[2]), .ZN(n367) );
  INV_X1 U190 ( .A(n369), .ZN(n368) );
  INV_X1 U191 ( .A(A[2]), .ZN(n377) );
  INV_X1 U192 ( .A(A[14]), .ZN(n381) );
  INV_X1 U193 ( .A(A[15]), .ZN(n382) );
  INV_X1 U194 ( .A(A[16]), .ZN(n383) );
  INV_X1 U195 ( .A(A[17]), .ZN(n384) );
  INV_X1 U196 ( .A(A[19]), .ZN(n385) );
  INV_X1 U197 ( .A(A[20]), .ZN(n386) );
  INV_X1 U198 ( .A(A[21]), .ZN(n387) );
  INV_X1 U199 ( .A(A[23]), .ZN(n388) );
  INV_X1 U200 ( .A(A[24]), .ZN(n389) );
  INV_X1 U201 ( .A(A[25]), .ZN(n390) );
  INV_X1 U202 ( .A(A[26]), .ZN(n391) );
  INV_X1 U203 ( .A(A[27]), .ZN(n392) );
  INV_X1 U204 ( .A(A[28]), .ZN(n393) );
  INV_X1 U205 ( .A(A[29]), .ZN(n394) );
  INV_X1 U206 ( .A(A[30]), .ZN(n395) );
  INV_X1 U207 ( .A(A[31]), .ZN(n396) );
endmodule


module SHIFTER_GENERIC_N32_DW_sla_0 ( A, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input SH_TC;
  wire   \A[0] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n22, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n111, n112, n113, n114, n116,
         n117, n118, n120, n121, n123, n126, n128, n129, n130, n131, n132,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n145, n147,
         n150, n151, n152, n155, n157, n159, n160, n161, n162, n164, n166,
         n167, n168, n170, n171, n172, n185, n288, n289, n324, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361;
  assign B[0] = \A[0] ;
  assign \A[0]  = A[0];

  NOR2_X2 U2 ( .A1(n336), .A2(SH[3]), .ZN(n73) );
  NOR2_X2 U3 ( .A1(SH[2]), .A2(SH[3]), .ZN(n75) );
  MUX2_X1 U143 ( .A(A[1]), .B(\A[0] ), .S(n34), .Z(n79) );
  AND2_X1 U4 ( .A1(n131), .A2(SH[2]), .ZN(n14) );
  INV_X1 U5 ( .A(n343), .ZN(n339) );
  INV_X1 U6 ( .A(n11), .ZN(n58) );
  NAND2_X1 U7 ( .A1(n343), .A2(\A[0] ), .ZN(n3) );
  INV_X1 U8 ( .A(n34), .ZN(n26) );
  NAND2_X1 U9 ( .A1(n73), .A2(n339), .ZN(n11) );
  INV_X1 U10 ( .A(n55), .ZN(n16) );
  OAI21_X1 U11 ( .B1(n341), .B2(n9), .A(n3), .ZN(B[3]) );
  OAI21_X1 U12 ( .B1(n340), .B2(n8), .A(n3), .ZN(B[4]) );
  OAI21_X1 U13 ( .B1(n342), .B2(n7), .A(n3), .ZN(B[5]) );
  OAI21_X1 U14 ( .B1(n342), .B2(n6), .A(n3), .ZN(B[6]) );
  OAI21_X1 U15 ( .B1(n342), .B2(n5), .A(n3), .ZN(B[7]) );
  OAI21_X1 U16 ( .B1(n342), .B2(n4), .A(n3), .ZN(B[8]) );
  OAI21_X1 U17 ( .B1(n342), .B2(n2), .A(n3), .ZN(B[9]) );
  OAI21_X1 U18 ( .B1(n341), .B2(n63), .A(n3), .ZN(B[10]) );
  OAI21_X1 U19 ( .B1(n340), .B2(n56), .A(n3), .ZN(B[11]) );
  OAI21_X1 U20 ( .B1(n341), .B2(n48), .A(n3), .ZN(B[12]) );
  OAI21_X1 U21 ( .B1(n341), .B2(n41), .A(n3), .ZN(B[13]) );
  OAI21_X1 U22 ( .B1(n340), .B2(n28), .A(n3), .ZN(B[14]) );
  OAI21_X1 U23 ( .B1(n340), .B2(n12), .A(n3), .ZN(B[15]) );
  INV_X1 U24 ( .A(n106), .ZN(n43) );
  INV_X1 U25 ( .A(n100), .ZN(n30) );
  INV_X1 U26 ( .A(n93), .ZN(n15) );
  BUF_X1 U27 ( .A(n338), .Z(n343) );
  INV_X1 U28 ( .A(A[1]), .ZN(n185) );
  OAI21_X1 U29 ( .B1(n341), .B2(n116), .A(n3), .ZN(B[1]) );
  OAI21_X1 U30 ( .B1(n340), .B2(n39), .A(n3), .ZN(B[2]) );
  INV_X1 U31 ( .A(n107), .ZN(n88) );
  BUF_X1 U32 ( .A(n338), .Z(n342) );
  BUF_X1 U33 ( .A(n337), .Z(n341) );
  BUF_X1 U34 ( .A(n337), .Z(n340) );
  INV_X1 U35 ( .A(n20), .ZN(n37) );
  INV_X1 U36 ( .A(n22), .ZN(n38) );
  OAI222_X1 U37 ( .A1(n34), .A2(n346), .B1(n185), .B2(n33), .C1(n344), .C2(
        n329), .ZN(n101) );
  NAND2_X1 U38 ( .A1(n75), .A2(n339), .ZN(n55) );
  INV_X1 U39 ( .A(n33), .ZN(n25) );
  AOI221_X1 U40 ( .B1(n25), .B2(A[16]), .C1(n26), .C2(n354), .A(n126), .ZN(
        n106) );
  OAI22_X1 U41 ( .A1(n352), .A2(n20), .B1(n351), .B2(n22), .ZN(n126) );
  AOI221_X1 U42 ( .B1(n25), .B2(n354), .C1(n26), .C2(A[18]), .A(n121), .ZN(
        n100) );
  OAI22_X1 U43 ( .A1(n353), .A2(n20), .B1(n352), .B2(n22), .ZN(n121) );
  AOI221_X1 U44 ( .B1(n25), .B2(A[18]), .C1(n26), .C2(A[19]), .A(n118), .ZN(
        n93) );
  OAI22_X1 U45 ( .A1(n355), .A2(n20), .B1(n353), .B2(n22), .ZN(n118) );
  AOI221_X1 U46 ( .B1(n79), .B2(n73), .C1(n72), .C2(n75), .A(n88), .ZN(n7) );
  AOI221_X1 U47 ( .B1(n101), .B2(n73), .C1(n102), .C2(n75), .A(n88), .ZN(n6)
         );
  AOI221_X1 U48 ( .B1(n94), .B2(n73), .C1(n95), .C2(n75), .A(n88), .ZN(n5) );
  AOI221_X1 U49 ( .B1(n86), .B2(n73), .C1(n87), .C2(n75), .A(n88), .ZN(n4) );
  AOI221_X1 U50 ( .B1(n72), .B2(n73), .C1(n74), .C2(n75), .A(n76), .ZN(n2) );
  INV_X1 U51 ( .A(n77), .ZN(n76) );
  AOI21_X1 U52 ( .B1(n78), .B2(n79), .A(n80), .ZN(n77) );
  AOI221_X1 U53 ( .B1(n102), .B2(n73), .C1(n99), .C2(n75), .A(n167), .ZN(n63)
         );
  INV_X1 U54 ( .A(n168), .ZN(n167) );
  AOI21_X1 U55 ( .B1(n78), .B2(n101), .A(n80), .ZN(n168) );
  AOI221_X1 U56 ( .B1(n74), .B2(n73), .C1(n70), .C2(n75), .A(n141), .ZN(n41)
         );
  INV_X1 U57 ( .A(n142), .ZN(n141) );
  AOI22_X1 U58 ( .A1(n136), .A2(n79), .B1(n78), .B2(n72), .ZN(n142) );
  AOI221_X1 U59 ( .B1(n99), .B2(n73), .C1(n65), .C2(n75), .A(n138), .ZN(n28)
         );
  INV_X1 U60 ( .A(n139), .ZN(n138) );
  AOI22_X1 U61 ( .A1(n136), .A2(n101), .B1(n78), .B2(n102), .ZN(n139) );
  NAND2_X1 U62 ( .A1(n335), .A2(n329), .ZN(n34) );
  OAI221_X1 U63 ( .B1(n106), .B2(n55), .C1(n116), .C2(n339), .A(n123), .ZN(
        B[17]) );
  AOI222_X1 U64 ( .A1(n58), .A2(n70), .B1(n18), .B2(n74), .C1(n14), .C2(n72), 
        .ZN(n123) );
  OAI221_X1 U65 ( .B1(n100), .B2(n55), .C1(n39), .C2(n339), .A(n120), .ZN(
        B[18]) );
  AOI222_X1 U66 ( .A1(n58), .A2(n65), .B1(n18), .B2(n99), .C1(n14), .C2(n102), 
        .ZN(n120) );
  OAI221_X1 U67 ( .B1(n93), .B2(n55), .C1(n9), .C2(n339), .A(n117), .ZN(B[19])
         );
  AOI222_X1 U68 ( .A1(n58), .A2(n59), .B1(n18), .B2(n92), .C1(n14), .C2(n95), 
        .ZN(n117) );
  OAI221_X1 U69 ( .B1(n85), .B2(n55), .C1(n8), .C2(n339), .A(n111), .ZN(B[20])
         );
  AOI222_X1 U70 ( .A1(n58), .A2(n50), .B1(n18), .B2(n84), .C1(n14), .C2(n87), 
        .ZN(n111) );
  OAI221_X1 U71 ( .B1(n71), .B2(n55), .C1(n7), .C2(n339), .A(n105), .ZN(B[21])
         );
  AOI222_X1 U72 ( .A1(n58), .A2(n43), .B1(n18), .B2(n70), .C1(n14), .C2(n74), 
        .ZN(n105) );
  OAI221_X1 U73 ( .B1(n66), .B2(n55), .C1(n6), .C2(n339), .A(n98), .ZN(B[22])
         );
  AOI222_X1 U74 ( .A1(n58), .A2(n30), .B1(n18), .B2(n65), .C1(n14), .C2(n99), 
        .ZN(n98) );
  OAI221_X1 U75 ( .B1(n60), .B2(n55), .C1(n5), .C2(n339), .A(n91), .ZN(B[23])
         );
  AOI222_X1 U76 ( .A1(n58), .A2(n15), .B1(n18), .B2(n59), .C1(n14), .C2(n92), 
        .ZN(n91) );
  OAI221_X1 U77 ( .B1(n47), .B2(n55), .C1(n4), .C2(n339), .A(n83), .ZN(B[24])
         );
  AOI222_X1 U78 ( .A1(n58), .A2(n52), .B1(n18), .B2(n50), .C1(n14), .C2(n84), 
        .ZN(n83) );
  OAI221_X1 U79 ( .B1(n40), .B2(n55), .C1(n2), .C2(n339), .A(n69), .ZN(B[25])
         );
  AOI222_X1 U80 ( .A1(n58), .A2(n45), .B1(n18), .B2(n43), .C1(n14), .C2(n70), 
        .ZN(n69) );
  OAI221_X1 U81 ( .B1(n27), .B2(n55), .C1(n63), .C2(n339), .A(n64), .ZN(B[26])
         );
  AOI222_X1 U82 ( .A1(n58), .A2(n32), .B1(n18), .B2(n30), .C1(n14), .C2(n65), 
        .ZN(n64) );
  OAI221_X1 U83 ( .B1(n10), .B2(n55), .C1(n56), .C2(n339), .A(n57), .ZN(B[27])
         );
  AOI222_X1 U84 ( .A1(n58), .A2(n19), .B1(n18), .B2(n15), .C1(n14), .C2(n59), 
        .ZN(n57) );
  OAI221_X1 U85 ( .B1(n128), .B2(n11), .C1(n112), .C2(n55), .A(n129), .ZN(
        B[16]) );
  INV_X1 U86 ( .A(n84), .ZN(n128) );
  AOI221_X1 U87 ( .B1(n14), .B2(n86), .C1(n18), .C2(n87), .A(n130), .ZN(n129)
         );
  INV_X1 U88 ( .A(n3), .ZN(n130) );
  AOI21_X1 U89 ( .B1(n94), .B2(n75), .A(n113), .ZN(n9) );
  AOI21_X1 U90 ( .B1(n86), .B2(n75), .A(n113), .ZN(n8) );
  AOI221_X1 U91 ( .B1(n92), .B2(n73), .C1(n59), .C2(n75), .A(n134), .ZN(n12)
         );
  INV_X1 U92 ( .A(n135), .ZN(n134) );
  AOI22_X1 U93 ( .A1(n136), .A2(n94), .B1(n78), .B2(n95), .ZN(n135) );
  AOI221_X1 U94 ( .B1(n95), .B2(n73), .C1(n92), .C2(n75), .A(n160), .ZN(n56)
         );
  INV_X1 U95 ( .A(n161), .ZN(n160) );
  AOI21_X1 U96 ( .B1(n78), .B2(n94), .A(n80), .ZN(n161) );
  AOI221_X1 U97 ( .B1(n87), .B2(n73), .C1(n84), .C2(n75), .A(n151), .ZN(n48)
         );
  INV_X1 U98 ( .A(n152), .ZN(n151) );
  AOI21_X1 U99 ( .B1(n78), .B2(n86), .A(n80), .ZN(n152) );
  INV_X1 U100 ( .A(n112), .ZN(n50) );
  INV_X1 U101 ( .A(n66), .ZN(n32) );
  INV_X1 U102 ( .A(n85), .ZN(n52) );
  INV_X1 U103 ( .A(n60), .ZN(n19) );
  INV_X1 U104 ( .A(n71), .ZN(n45) );
  BUF_X1 U105 ( .A(SH[4]), .Z(n338) );
  OAI21_X1 U106 ( .B1(n344), .B2(n336), .A(n107), .ZN(n113) );
  NOR2_X1 U107 ( .A1(n336), .A2(n107), .ZN(n80) );
  AND2_X1 U108 ( .A1(n131), .A2(n336), .ZN(n18) );
  AND2_X1 U109 ( .A1(SH[3]), .A2(n336), .ZN(n78) );
  AOI21_X1 U110 ( .B1(n79), .B2(n75), .A(n113), .ZN(n116) );
  AOI21_X1 U111 ( .B1(n101), .B2(n75), .A(n113), .ZN(n39) );
  NAND2_X1 U112 ( .A1(SH[3]), .A2(\A[0] ), .ZN(n107) );
  INV_X1 U113 ( .A(n289), .ZN(n288) );
  AND2_X1 U114 ( .A1(SH[3]), .A2(n339), .ZN(n131) );
  BUF_X1 U115 ( .A(SH[4]), .Z(n337) );
  NAND2_X1 U116 ( .A1(SH[0]), .A2(n329), .ZN(n33) );
  OAI221_X1 U117 ( .B1(n33), .B2(n347), .C1(n34), .C2(n332), .A(n159), .ZN(n87) );
  AOI22_X1 U118 ( .A1(A[6]), .A2(n37), .B1(A[5]), .B2(n38), .ZN(n159) );
  OAI221_X1 U119 ( .B1(n33), .B2(n289), .C1(n34), .C2(n330), .A(n145), .ZN(n72) );
  AOI22_X1 U120 ( .A1(A[3]), .A2(n37), .B1(A[2]), .B2(n38), .ZN(n145) );
  OAI221_X1 U121 ( .B1(n33), .B2(n331), .C1(n34), .C2(n347), .A(n166), .ZN(n95) );
  AOI22_X1 U122 ( .A1(A[5]), .A2(n37), .B1(n288), .B2(n38), .ZN(n166) );
  OAI221_X1 U123 ( .B1(n33), .B2(n348), .C1(n34), .C2(n349), .A(n170), .ZN(n99) );
  AOI22_X1 U124 ( .A1(A[8]), .A2(n37), .B1(A[7]), .B2(n38), .ZN(n170) );
  OAI221_X1 U125 ( .B1(n33), .B2(n350), .C1(n34), .C2(n351), .A(n140), .ZN(n65) );
  AOI22_X1 U126 ( .A1(A[12]), .A2(n37), .B1(A[11]), .B2(n38), .ZN(n140) );
  OAI221_X1 U127 ( .B1(n33), .B2(n351), .C1(n34), .C2(n352), .A(n137), .ZN(n59) );
  AOI22_X1 U128 ( .A1(A[13]), .A2(n37), .B1(A[12]), .B2(n38), .ZN(n137) );
  OAI221_X1 U129 ( .B1(n185), .B2(n20), .C1(n345), .C2(n22), .A(n162), .ZN(n94) );
  AOI22_X1 U130 ( .A1(n25), .A2(A[2]), .B1(A[3]), .B2(n26), .ZN(n162) );
  OAI221_X1 U131 ( .B1(n20), .B2(n346), .C1(n185), .C2(n22), .A(n155), .ZN(n86) );
  AOI22_X1 U132 ( .A1(n25), .A2(A[3]), .B1(n288), .B2(n26), .ZN(n155) );
  AOI221_X1 U133 ( .B1(n25), .B2(A[24]), .C1(n26), .C2(A[25]), .A(n81), .ZN(
        n40) );
  INV_X1 U134 ( .A(n82), .ZN(n81) );
  AOI22_X1 U135 ( .A1(A[23]), .A2(n37), .B1(A[22]), .B2(n38), .ZN(n82) );
  AOI221_X1 U136 ( .B1(n25), .B2(A[21]), .C1(n26), .C2(A[22]), .A(n103), .ZN(
        n66) );
  INV_X1 U137 ( .A(n104), .ZN(n103) );
  AOI22_X1 U138 ( .A1(A[20]), .A2(n37), .B1(A[19]), .B2(n38), .ZN(n104) );
  AOI221_X1 U139 ( .B1(n25), .B2(A[19]), .C1(n26), .C2(A[20]), .A(n114), .ZN(
        n85) );
  OAI22_X1 U140 ( .A1(n324), .A2(n20), .B1(n355), .B2(n22), .ZN(n114) );
  AOI221_X1 U141 ( .B1(n25), .B2(A[22]), .C1(n26), .C2(A[23]), .A(n96), .ZN(
        n60) );
  INV_X1 U142 ( .A(n97), .ZN(n96) );
  AOI22_X1 U144 ( .A1(A[21]), .A2(n37), .B1(A[20]), .B2(n38), .ZN(n97) );
  AOI221_X1 U145 ( .B1(n25), .B2(A[20]), .C1(n26), .C2(A[21]), .A(n108), .ZN(
        n71) );
  OAI22_X1 U146 ( .A1(n356), .A2(n20), .B1(n324), .B2(n22), .ZN(n108) );
  AOI221_X1 U147 ( .B1(n25), .B2(A[15]), .C1(n26), .C2(A[16]), .A(n132), .ZN(
        n112) );
  OAI22_X1 U148 ( .A1(n351), .A2(n20), .B1(n350), .B2(n22), .ZN(n132) );
  NAND2_X1 U149 ( .A1(SH[1]), .A2(n335), .ZN(n20) );
  NAND2_X1 U150 ( .A1(SH[0]), .A2(SH[1]), .ZN(n22) );
  INV_X1 U151 ( .A(n171), .ZN(n102) );
  AOI221_X1 U152 ( .B1(n37), .B2(n288), .C1(A[3]), .C2(n38), .A(n172), .ZN(
        n171) );
  OAI22_X1 U153 ( .A1(n330), .A2(n33), .B1(n331), .B2(n34), .ZN(n172) );
  OAI221_X1 U154 ( .B1(n47), .B2(n11), .C1(n48), .C2(n339), .A(n49), .ZN(B[28]) );
  AOI222_X1 U155 ( .A1(n14), .A2(n50), .B1(n16), .B2(n51), .C1(n18), .C2(n52), 
        .ZN(n49) );
  OAI221_X1 U156 ( .B1(n33), .B2(n358), .C1(n34), .C2(n359), .A(n54), .ZN(n51)
         );
  AOI22_X1 U157 ( .A1(A[26]), .A2(n37), .B1(A[25]), .B2(n38), .ZN(n54) );
  OAI221_X1 U158 ( .B1(n40), .B2(n11), .C1(n41), .C2(n339), .A(n42), .ZN(B[29]) );
  AOI222_X1 U159 ( .A1(n14), .A2(n43), .B1(n16), .B2(n44), .C1(n18), .C2(n45), 
        .ZN(n42) );
  OAI221_X1 U160 ( .B1(n33), .B2(n359), .C1(n34), .C2(n360), .A(n46), .ZN(n44)
         );
  AOI22_X1 U161 ( .A1(n357), .A2(n37), .B1(A[26]), .B2(n38), .ZN(n46) );
  OAI221_X1 U162 ( .B1(n27), .B2(n11), .C1(n28), .C2(n339), .A(n29), .ZN(B[30]) );
  AOI222_X1 U163 ( .A1(n14), .A2(n30), .B1(n16), .B2(n31), .C1(n18), .C2(n32), 
        .ZN(n29) );
  OAI221_X1 U164 ( .B1(n33), .B2(n360), .C1(n34), .C2(n361), .A(n36), .ZN(n31)
         );
  OAI221_X1 U165 ( .B1(n10), .B2(n11), .C1(n12), .C2(n339), .A(n13), .ZN(B[31]) );
  AOI222_X1 U166 ( .A1(n14), .A2(n15), .B1(n16), .B2(n17), .C1(n18), .C2(n19), 
        .ZN(n13) );
  OAI221_X1 U167 ( .B1(n20), .B2(n360), .C1(n22), .C2(n359), .A(n24), .ZN(n17)
         );
  AOI22_X1 U168 ( .A1(A[30]), .A2(n25), .B1(A[31]), .B2(n26), .ZN(n24) );
  AOI221_X1 U169 ( .B1(n25), .B2(A[23]), .C1(n26), .C2(A[24]), .A(n89), .ZN(
        n47) );
  INV_X1 U170 ( .A(n90), .ZN(n89) );
  AOI22_X1 U171 ( .A1(A[22]), .A2(n37), .B1(A[21]), .B2(n38), .ZN(n90) );
  AOI22_X1 U172 ( .A1(A[28]), .A2(n37), .B1(n357), .B2(n38), .ZN(n36) );
  OAI221_X1 U173 ( .B1(n33), .B2(n333), .C1(n34), .C2(n334), .A(n157), .ZN(n84) );
  AOI22_X1 U174 ( .A1(A[10]), .A2(n37), .B1(A[9]), .B2(n38), .ZN(n157) );
  OAI221_X1 U175 ( .B1(n33), .B2(n334), .C1(n34), .C2(n350), .A(n147), .ZN(n70) );
  AOI22_X1 U176 ( .A1(A[11]), .A2(n37), .B1(A[10]), .B2(n38), .ZN(n147) );
  OAI221_X1 U177 ( .B1(n33), .B2(n332), .C1(n34), .C2(n348), .A(n150), .ZN(n74) );
  AOI22_X1 U178 ( .A1(A[7]), .A2(n37), .B1(A[6]), .B2(n38), .ZN(n150) );
  OAI221_X1 U179 ( .B1(n33), .B2(n349), .C1(n34), .C2(n333), .A(n164), .ZN(n92) );
  AOI22_X1 U180 ( .A1(A[9]), .A2(n37), .B1(A[8]), .B2(n38), .ZN(n164) );
  AOI221_X1 U181 ( .B1(n25), .B2(A[26]), .C1(n26), .C2(n357), .A(n61), .ZN(n10) );
  INV_X1 U182 ( .A(n62), .ZN(n61) );
  AOI22_X1 U183 ( .A1(A[25]), .A2(n37), .B1(A[24]), .B2(n38), .ZN(n62) );
  AOI221_X1 U184 ( .B1(n25), .B2(A[25]), .C1(n26), .C2(A[26]), .A(n67), .ZN(
        n27) );
  INV_X1 U185 ( .A(n68), .ZN(n67) );
  AOI22_X1 U186 ( .A1(A[24]), .A2(n37), .B1(A[23]), .B2(n38), .ZN(n68) );
  INV_X1 U187 ( .A(A[16]), .ZN(n353) );
  INV_X1 U188 ( .A(A[17]), .ZN(n355) );
  INV_X1 U189 ( .A(A[18]), .ZN(n324) );
  INV_X1 U190 ( .A(A[4]), .ZN(n289) );
  AND2_X1 U191 ( .A1(SH[2]), .A2(SH[3]), .ZN(n136) );
  INV_X1 U192 ( .A(SH[1]), .ZN(n329) );
  INV_X1 U193 ( .A(A[5]), .ZN(n330) );
  INV_X1 U194 ( .A(A[6]), .ZN(n331) );
  INV_X1 U195 ( .A(A[8]), .ZN(n332) );
  INV_X1 U196 ( .A(A[11]), .ZN(n333) );
  INV_X1 U197 ( .A(A[12]), .ZN(n334) );
  INV_X1 U198 ( .A(A[2]), .ZN(n346) );
  INV_X1 U199 ( .A(SH[0]), .ZN(n335) );
  INV_X1 U200 ( .A(SH[2]), .ZN(n336) );
  INV_X1 U201 ( .A(\A[0] ), .ZN(n344) );
  INV_X1 U202 ( .A(\A[0] ), .ZN(n345) );
  INV_X1 U203 ( .A(A[7]), .ZN(n347) );
  INV_X1 U204 ( .A(A[9]), .ZN(n348) );
  INV_X1 U205 ( .A(A[10]), .ZN(n349) );
  INV_X1 U206 ( .A(A[13]), .ZN(n350) );
  INV_X1 U207 ( .A(A[14]), .ZN(n351) );
  INV_X1 U208 ( .A(A[15]), .ZN(n352) );
  INV_X1 U209 ( .A(n355), .ZN(n354) );
  INV_X1 U210 ( .A(A[19]), .ZN(n356) );
  INV_X1 U211 ( .A(n358), .ZN(n357) );
  INV_X1 U212 ( .A(A[27]), .ZN(n358) );
  INV_X1 U213 ( .A(A[28]), .ZN(n359) );
  INV_X1 U214 ( .A(A[29]), .ZN(n360) );
  INV_X1 U215 ( .A(A[30]), .ZN(n361) );
endmodule


module SHIFTER_GENERIC_N32_DW01_ash_0 ( A, DATA_TC, SH, SH_TC, B );
  input [31:0] A;
  input [4:0] SH;
  output [31:0] B;
  input DATA_TC, SH_TC;
  wire   \ML_int[1][31] , \ML_int[1][30] , \ML_int[1][29] , \ML_int[1][28] ,
         \ML_int[1][27] , \ML_int[1][26] , \ML_int[1][25] , \ML_int[1][24] ,
         \ML_int[1][23] , \ML_int[1][22] , \ML_int[1][21] , \ML_int[1][20] ,
         \ML_int[1][19] , \ML_int[1][18] , \ML_int[1][17] , \ML_int[1][16] ,
         \ML_int[1][15] , \ML_int[1][14] , \ML_int[1][13] , \ML_int[1][12] ,
         \ML_int[1][11] , \ML_int[1][10] , \ML_int[1][9] , \ML_int[1][8] ,
         \ML_int[1][7] , \ML_int[1][6] , \ML_int[1][5] , \ML_int[1][4] ,
         \ML_int[1][3] , \ML_int[1][2] , \ML_int[1][1] , \ML_int[1][0] ,
         \ML_int[2][31] , \ML_int[2][30] , \ML_int[2][29] , \ML_int[2][28] ,
         \ML_int[2][27] , \ML_int[2][26] , \ML_int[2][25] , \ML_int[2][24] ,
         \ML_int[2][23] , \ML_int[2][22] , \ML_int[2][21] , \ML_int[2][20] ,
         \ML_int[2][19] , \ML_int[2][18] , \ML_int[2][17] , \ML_int[2][16] ,
         \ML_int[2][15] , \ML_int[2][14] , \ML_int[2][13] , \ML_int[2][12] ,
         \ML_int[2][11] , \ML_int[2][10] , \ML_int[2][9] , \ML_int[2][8] ,
         \ML_int[2][7] , \ML_int[2][6] , \ML_int[2][5] , \ML_int[2][4] ,
         \ML_int[2][3] , \ML_int[2][2] , \ML_int[2][1] , \ML_int[2][0] ,
         \ML_int[3][31] , \ML_int[3][30] , \ML_int[3][29] , \ML_int[3][28] ,
         \ML_int[3][27] , \ML_int[3][26] , \ML_int[3][25] , \ML_int[3][24] ,
         \ML_int[3][23] , \ML_int[3][22] , \ML_int[3][21] , \ML_int[3][20] ,
         \ML_int[3][19] , \ML_int[3][18] , \ML_int[3][17] , \ML_int[3][16] ,
         \ML_int[3][15] , \ML_int[3][14] , \ML_int[3][13] , \ML_int[3][12] ,
         \ML_int[3][11] , \ML_int[3][10] , \ML_int[3][9] , \ML_int[3][8] ,
         \ML_int[3][7] , \ML_int[3][6] , \ML_int[3][5] , \ML_int[3][4] ,
         \ML_int[3][3] , \ML_int[3][2] , \ML_int[3][1] , \ML_int[3][0] ,
         \ML_int[4][31] , \ML_int[4][30] , \ML_int[4][29] , \ML_int[4][28] ,
         \ML_int[4][27] , \ML_int[4][26] , \ML_int[4][25] , \ML_int[4][24] ,
         \ML_int[4][23] , \ML_int[4][22] , \ML_int[4][21] , \ML_int[4][20] ,
         \ML_int[4][19] , \ML_int[4][18] , \ML_int[4][17] , \ML_int[4][16] ,
         \ML_int[4][15] , \ML_int[4][14] , \ML_int[4][13] , \ML_int[4][12] ,
         \ML_int[4][11] , \ML_int[4][10] , \ML_int[4][9] , \ML_int[4][8] ,
         \ML_int[4][7] , \ML_int[4][6] , \ML_int[4][5] , \ML_int[4][4] ,
         \ML_int[4][3] , \ML_int[4][2] , \ML_int[4][1] , \ML_int[4][0] , n3,
         n4, n5, n6, n7, n8, n9, n10, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87;

  MUX2_X1 M1_4_31 ( .A(\ML_int[4][31] ), .B(\ML_int[4][15] ), .S(SH[4]), .Z(
        B[31]) );
  MUX2_X1 M1_4_30 ( .A(\ML_int[4][30] ), .B(\ML_int[4][14] ), .S(SH[4]), .Z(
        B[30]) );
  MUX2_X1 M1_4_29 ( .A(\ML_int[4][29] ), .B(\ML_int[4][13] ), .S(SH[4]), .Z(
        B[29]) );
  MUX2_X1 M1_4_28 ( .A(\ML_int[4][28] ), .B(\ML_int[4][12] ), .S(SH[4]), .Z(
        B[28]) );
  MUX2_X1 M1_4_27 ( .A(\ML_int[4][27] ), .B(\ML_int[4][11] ), .S(SH[4]), .Z(
        B[27]) );
  MUX2_X1 M1_4_26 ( .A(\ML_int[4][26] ), .B(\ML_int[4][10] ), .S(SH[4]), .Z(
        B[26]) );
  MUX2_X1 M1_4_25 ( .A(\ML_int[4][25] ), .B(\ML_int[4][9] ), .S(SH[4]), .Z(
        B[25]) );
  MUX2_X1 M1_4_24 ( .A(\ML_int[4][24] ), .B(\ML_int[4][8] ), .S(n86), .Z(B[24]) );
  MUX2_X1 M1_4_23 ( .A(\ML_int[4][23] ), .B(\ML_int[4][7] ), .S(SH[4]), .Z(
        B[23]) );
  MUX2_X1 M1_4_22 ( .A(\ML_int[4][22] ), .B(\ML_int[4][6] ), .S(n86), .Z(B[22]) );
  MUX2_X1 M1_4_21 ( .A(\ML_int[4][21] ), .B(\ML_int[4][5] ), .S(n86), .Z(B[21]) );
  MUX2_X1 M1_4_20 ( .A(\ML_int[4][20] ), .B(\ML_int[4][4] ), .S(n86), .Z(B[20]) );
  MUX2_X1 M1_4_19 ( .A(\ML_int[4][19] ), .B(\ML_int[4][3] ), .S(SH[4]), .Z(
        B[19]) );
  MUX2_X1 M1_4_18 ( .A(\ML_int[4][18] ), .B(\ML_int[4][2] ), .S(n86), .Z(B[18]) );
  MUX2_X1 M1_4_17 ( .A(\ML_int[4][17] ), .B(\ML_int[4][1] ), .S(SH[4]), .Z(
        B[17]) );
  MUX2_X1 M1_4_16 ( .A(\ML_int[4][16] ), .B(\ML_int[4][0] ), .S(SH[4]), .Z(
        B[16]) );
  MUX2_X1 M1_3_31 ( .A(\ML_int[3][31] ), .B(\ML_int[3][23] ), .S(n84), .Z(
        \ML_int[4][31] ) );
  MUX2_X1 M1_3_30 ( .A(\ML_int[3][30] ), .B(\ML_int[3][22] ), .S(n84), .Z(
        \ML_int[4][30] ) );
  MUX2_X1 M1_3_29 ( .A(\ML_int[3][29] ), .B(\ML_int[3][21] ), .S(n83), .Z(
        \ML_int[4][29] ) );
  MUX2_X1 M1_3_28 ( .A(\ML_int[3][28] ), .B(\ML_int[3][20] ), .S(n83), .Z(
        \ML_int[4][28] ) );
  MUX2_X1 M1_3_27 ( .A(\ML_int[3][27] ), .B(\ML_int[3][19] ), .S(n83), .Z(
        \ML_int[4][27] ) );
  MUX2_X1 M1_3_26 ( .A(\ML_int[3][26] ), .B(\ML_int[3][18] ), .S(n83), .Z(
        \ML_int[4][26] ) );
  MUX2_X1 M1_3_25 ( .A(\ML_int[3][25] ), .B(\ML_int[3][17] ), .S(n83), .Z(
        \ML_int[4][25] ) );
  MUX2_X1 M1_3_24 ( .A(\ML_int[3][24] ), .B(\ML_int[3][16] ), .S(n83), .Z(
        \ML_int[4][24] ) );
  MUX2_X1 M1_3_23 ( .A(\ML_int[3][23] ), .B(\ML_int[3][15] ), .S(n83), .Z(
        \ML_int[4][23] ) );
  MUX2_X1 M1_3_22 ( .A(\ML_int[3][22] ), .B(\ML_int[3][14] ), .S(n83), .Z(
        \ML_int[4][22] ) );
  MUX2_X1 M1_3_21 ( .A(\ML_int[3][21] ), .B(\ML_int[3][13] ), .S(n83), .Z(
        \ML_int[4][21] ) );
  MUX2_X1 M1_3_20 ( .A(\ML_int[3][20] ), .B(\ML_int[3][12] ), .S(n83), .Z(
        \ML_int[4][20] ) );
  MUX2_X1 M1_3_19 ( .A(\ML_int[3][19] ), .B(\ML_int[3][11] ), .S(n84), .Z(
        \ML_int[4][19] ) );
  MUX2_X1 M1_3_18 ( .A(\ML_int[3][18] ), .B(\ML_int[3][10] ), .S(SH[3]), .Z(
        \ML_int[4][18] ) );
  MUX2_X1 M1_3_17 ( .A(\ML_int[3][17] ), .B(\ML_int[3][9] ), .S(n83), .Z(
        \ML_int[4][17] ) );
  MUX2_X1 M1_3_16 ( .A(\ML_int[3][16] ), .B(\ML_int[3][8] ), .S(n84), .Z(
        \ML_int[4][16] ) );
  MUX2_X1 M1_3_15 ( .A(\ML_int[3][15] ), .B(\ML_int[3][7] ), .S(n84), .Z(
        \ML_int[4][15] ) );
  MUX2_X1 M1_3_14 ( .A(\ML_int[3][14] ), .B(\ML_int[3][6] ), .S(n84), .Z(
        \ML_int[4][14] ) );
  MUX2_X1 M1_3_13 ( .A(\ML_int[3][13] ), .B(\ML_int[3][5] ), .S(n84), .Z(
        \ML_int[4][13] ) );
  MUX2_X1 M1_3_12 ( .A(\ML_int[3][12] ), .B(\ML_int[3][4] ), .S(n84), .Z(
        \ML_int[4][12] ) );
  MUX2_X1 M1_3_11 ( .A(\ML_int[3][11] ), .B(\ML_int[3][3] ), .S(n84), .Z(
        \ML_int[4][11] ) );
  MUX2_X1 M1_3_10 ( .A(\ML_int[3][10] ), .B(\ML_int[3][2] ), .S(n84), .Z(
        \ML_int[4][10] ) );
  MUX2_X1 M1_3_9 ( .A(\ML_int[3][9] ), .B(\ML_int[3][1] ), .S(n84), .Z(
        \ML_int[4][9] ) );
  MUX2_X1 M1_3_8 ( .A(\ML_int[3][8] ), .B(\ML_int[3][0] ), .S(n83), .Z(
        \ML_int[4][8] ) );
  MUX2_X1 M1_2_31 ( .A(\ML_int[2][31] ), .B(\ML_int[2][27] ), .S(SH[2]), .Z(
        \ML_int[3][31] ) );
  MUX2_X1 M1_2_30 ( .A(\ML_int[2][30] ), .B(\ML_int[2][26] ), .S(SH[2]), .Z(
        \ML_int[3][30] ) );
  MUX2_X1 M1_2_29 ( .A(\ML_int[2][29] ), .B(\ML_int[2][25] ), .S(n80), .Z(
        \ML_int[3][29] ) );
  MUX2_X1 M1_2_28 ( .A(\ML_int[2][28] ), .B(\ML_int[2][24] ), .S(n81), .Z(
        \ML_int[3][28] ) );
  MUX2_X1 M1_2_27 ( .A(\ML_int[2][27] ), .B(\ML_int[2][23] ), .S(SH[2]), .Z(
        \ML_int[3][27] ) );
  MUX2_X1 M1_2_26 ( .A(\ML_int[2][26] ), .B(\ML_int[2][22] ), .S(n81), .Z(
        \ML_int[3][26] ) );
  MUX2_X1 M1_2_25 ( .A(\ML_int[2][25] ), .B(\ML_int[2][21] ), .S(n81), .Z(
        \ML_int[3][25] ) );
  MUX2_X1 M1_2_24 ( .A(\ML_int[2][24] ), .B(\ML_int[2][20] ), .S(n81), .Z(
        \ML_int[3][24] ) );
  MUX2_X1 M1_2_23 ( .A(\ML_int[2][23] ), .B(\ML_int[2][19] ), .S(n81), .Z(
        \ML_int[3][23] ) );
  MUX2_X1 M1_2_22 ( .A(\ML_int[2][22] ), .B(\ML_int[2][18] ), .S(n81), .Z(
        \ML_int[3][22] ) );
  MUX2_X1 M1_2_21 ( .A(\ML_int[2][21] ), .B(\ML_int[2][17] ), .S(n81), .Z(
        \ML_int[3][21] ) );
  MUX2_X1 M1_2_20 ( .A(\ML_int[2][20] ), .B(\ML_int[2][16] ), .S(n81), .Z(
        \ML_int[3][20] ) );
  MUX2_X1 M1_2_19 ( .A(\ML_int[2][19] ), .B(\ML_int[2][15] ), .S(n81), .Z(
        \ML_int[3][19] ) );
  MUX2_X1 M1_2_18 ( .A(\ML_int[2][18] ), .B(\ML_int[2][14] ), .S(n81), .Z(
        \ML_int[3][18] ) );
  MUX2_X1 M1_2_17 ( .A(\ML_int[2][17] ), .B(\ML_int[2][13] ), .S(SH[2]), .Z(
        \ML_int[3][17] ) );
  MUX2_X1 M1_2_16 ( .A(\ML_int[2][16] ), .B(\ML_int[2][12] ), .S(SH[2]), .Z(
        \ML_int[3][16] ) );
  MUX2_X1 M1_2_15 ( .A(\ML_int[2][15] ), .B(\ML_int[2][11] ), .S(SH[2]), .Z(
        \ML_int[3][15] ) );
  MUX2_X1 M1_2_14 ( .A(\ML_int[2][14] ), .B(\ML_int[2][10] ), .S(n80), .Z(
        \ML_int[3][14] ) );
  MUX2_X1 M1_2_13 ( .A(\ML_int[2][13] ), .B(\ML_int[2][9] ), .S(n80), .Z(
        \ML_int[3][13] ) );
  MUX2_X1 M1_2_12 ( .A(\ML_int[2][12] ), .B(\ML_int[2][8] ), .S(n80), .Z(
        \ML_int[3][12] ) );
  MUX2_X1 M1_2_11 ( .A(\ML_int[2][11] ), .B(\ML_int[2][7] ), .S(n80), .Z(
        \ML_int[3][11] ) );
  MUX2_X1 M1_2_10 ( .A(\ML_int[2][10] ), .B(\ML_int[2][6] ), .S(n80), .Z(
        \ML_int[3][10] ) );
  MUX2_X1 M1_2_9 ( .A(\ML_int[2][9] ), .B(\ML_int[2][5] ), .S(n80), .Z(
        \ML_int[3][9] ) );
  MUX2_X1 M1_2_8 ( .A(\ML_int[2][8] ), .B(\ML_int[2][4] ), .S(n80), .Z(
        \ML_int[3][8] ) );
  MUX2_X1 M1_2_7 ( .A(\ML_int[2][7] ), .B(\ML_int[2][3] ), .S(n80), .Z(
        \ML_int[3][7] ) );
  MUX2_X1 M1_2_6 ( .A(\ML_int[2][6] ), .B(\ML_int[2][2] ), .S(n80), .Z(
        \ML_int[3][6] ) );
  MUX2_X1 M1_2_5 ( .A(\ML_int[2][5] ), .B(\ML_int[2][1] ), .S(n80), .Z(
        \ML_int[3][5] ) );
  MUX2_X1 M1_2_4 ( .A(\ML_int[2][4] ), .B(\ML_int[2][0] ), .S(n81), .Z(
        \ML_int[3][4] ) );
  MUX2_X1 M1_1_31 ( .A(\ML_int[1][31] ), .B(\ML_int[1][29] ), .S(n74), .Z(
        \ML_int[2][31] ) );
  MUX2_X1 M1_1_30 ( .A(\ML_int[1][30] ), .B(\ML_int[1][28] ), .S(n75), .Z(
        \ML_int[2][30] ) );
  MUX2_X1 M1_1_29 ( .A(\ML_int[1][29] ), .B(\ML_int[1][27] ), .S(n75), .Z(
        \ML_int[2][29] ) );
  MUX2_X1 M1_1_28 ( .A(\ML_int[1][28] ), .B(\ML_int[1][26] ), .S(n74), .Z(
        \ML_int[2][28] ) );
  MUX2_X1 M1_1_27 ( .A(\ML_int[1][27] ), .B(\ML_int[1][25] ), .S(SH[1]), .Z(
        \ML_int[2][27] ) );
  MUX2_X1 M1_1_26 ( .A(\ML_int[1][26] ), .B(\ML_int[1][24] ), .S(SH[1]), .Z(
        \ML_int[2][26] ) );
  MUX2_X1 M1_1_25 ( .A(\ML_int[1][25] ), .B(\ML_int[1][23] ), .S(SH[1]), .Z(
        \ML_int[2][25] ) );
  MUX2_X1 M1_1_24 ( .A(\ML_int[1][24] ), .B(\ML_int[1][22] ), .S(n75), .Z(
        \ML_int[2][24] ) );
  MUX2_X1 M1_1_23 ( .A(\ML_int[1][23] ), .B(\ML_int[1][21] ), .S(n75), .Z(
        \ML_int[2][23] ) );
  MUX2_X1 M1_1_22 ( .A(\ML_int[1][22] ), .B(\ML_int[1][20] ), .S(n75), .Z(
        \ML_int[2][22] ) );
  MUX2_X1 M1_1_21 ( .A(\ML_int[1][21] ), .B(\ML_int[1][19] ), .S(n75), .Z(
        \ML_int[2][21] ) );
  MUX2_X1 M1_1_20 ( .A(\ML_int[1][20] ), .B(\ML_int[1][18] ), .S(n75), .Z(
        \ML_int[2][20] ) );
  MUX2_X1 M1_1_19 ( .A(\ML_int[1][19] ), .B(\ML_int[1][17] ), .S(n75), .Z(
        \ML_int[2][19] ) );
  MUX2_X1 M1_1_18 ( .A(\ML_int[1][18] ), .B(\ML_int[1][16] ), .S(n75), .Z(
        \ML_int[2][18] ) );
  MUX2_X1 M1_1_17 ( .A(\ML_int[1][17] ), .B(\ML_int[1][15] ), .S(n75), .Z(
        \ML_int[2][17] ) );
  MUX2_X1 M1_1_16 ( .A(\ML_int[1][16] ), .B(\ML_int[1][14] ), .S(n74), .Z(
        \ML_int[2][16] ) );
  MUX2_X1 M1_1_15 ( .A(\ML_int[1][15] ), .B(\ML_int[1][13] ), .S(n75), .Z(
        \ML_int[2][15] ) );
  MUX2_X1 M1_1_14 ( .A(\ML_int[1][14] ), .B(\ML_int[1][12] ), .S(n74), .Z(
        \ML_int[2][14] ) );
  MUX2_X1 M1_1_13 ( .A(\ML_int[1][13] ), .B(\ML_int[1][11] ), .S(SH[1]), .Z(
        \ML_int[2][13] ) );
  MUX2_X1 M1_1_12 ( .A(\ML_int[1][12] ), .B(\ML_int[1][10] ), .S(n74), .Z(
        \ML_int[2][12] ) );
  MUX2_X1 M1_1_11 ( .A(\ML_int[1][11] ), .B(\ML_int[1][9] ), .S(n74), .Z(
        \ML_int[2][11] ) );
  MUX2_X1 M1_1_10 ( .A(\ML_int[1][10] ), .B(\ML_int[1][8] ), .S(n74), .Z(
        \ML_int[2][10] ) );
  MUX2_X1 M1_1_9 ( .A(\ML_int[1][9] ), .B(\ML_int[1][7] ), .S(n74), .Z(
        \ML_int[2][9] ) );
  MUX2_X1 M1_1_8 ( .A(\ML_int[1][8] ), .B(\ML_int[1][6] ), .S(n74), .Z(
        \ML_int[2][8] ) );
  MUX2_X1 M1_1_7 ( .A(\ML_int[1][7] ), .B(\ML_int[1][5] ), .S(n74), .Z(
        \ML_int[2][7] ) );
  MUX2_X1 M1_1_6 ( .A(\ML_int[1][6] ), .B(\ML_int[1][4] ), .S(n74), .Z(
        \ML_int[2][6] ) );
  MUX2_X1 M1_1_5 ( .A(\ML_int[1][5] ), .B(\ML_int[1][3] ), .S(n74), .Z(
        \ML_int[2][5] ) );
  MUX2_X1 M1_1_4 ( .A(\ML_int[1][4] ), .B(\ML_int[1][2] ), .S(n74), .Z(
        \ML_int[2][4] ) );
  MUX2_X1 M1_1_3 ( .A(\ML_int[1][3] ), .B(\ML_int[1][1] ), .S(n75), .Z(
        \ML_int[2][3] ) );
  MUX2_X1 M1_1_2 ( .A(\ML_int[1][2] ), .B(\ML_int[1][0] ), .S(n75), .Z(
        \ML_int[2][2] ) );
  MUX2_X1 M1_0_31 ( .A(A[31]), .B(A[30]), .S(SH[0]), .Z(\ML_int[1][31] ) );
  MUX2_X1 M1_0_30 ( .A(A[30]), .B(A[29]), .S(SH[0]), .Z(\ML_int[1][30] ) );
  MUX2_X1 M1_0_29 ( .A(A[29]), .B(A[28]), .S(n78), .Z(\ML_int[1][29] ) );
  MUX2_X1 M1_0_28 ( .A(A[28]), .B(A[27]), .S(n78), .Z(\ML_int[1][28] ) );
  MUX2_X1 M1_0_27 ( .A(A[27]), .B(A[26]), .S(n78), .Z(\ML_int[1][27] ) );
  MUX2_X1 M1_0_26 ( .A(A[26]), .B(A[25]), .S(n78), .Z(\ML_int[1][26] ) );
  MUX2_X1 M1_0_25 ( .A(A[25]), .B(A[24]), .S(n78), .Z(\ML_int[1][25] ) );
  MUX2_X1 M1_0_24 ( .A(A[24]), .B(A[23]), .S(n78), .Z(\ML_int[1][24] ) );
  MUX2_X1 M1_0_23 ( .A(A[23]), .B(A[22]), .S(n78), .Z(\ML_int[1][23] ) );
  MUX2_X1 M1_0_22 ( .A(A[22]), .B(A[21]), .S(n77), .Z(\ML_int[1][22] ) );
  MUX2_X1 M1_0_21 ( .A(A[21]), .B(A[20]), .S(SH[0]), .Z(\ML_int[1][21] ) );
  MUX2_X1 M1_0_20 ( .A(A[20]), .B(A[19]), .S(SH[0]), .Z(\ML_int[1][20] ) );
  MUX2_X1 M1_0_19 ( .A(A[19]), .B(A[18]), .S(SH[0]), .Z(\ML_int[1][19] ) );
  MUX2_X1 M1_0_18 ( .A(A[18]), .B(A[17]), .S(SH[0]), .Z(\ML_int[1][18] ) );
  MUX2_X1 M1_0_17 ( .A(A[17]), .B(A[16]), .S(n78), .Z(\ML_int[1][17] ) );
  MUX2_X1 M1_0_16 ( .A(A[16]), .B(A[15]), .S(SH[0]), .Z(\ML_int[1][16] ) );
  MUX2_X1 M1_0_15 ( .A(A[15]), .B(A[14]), .S(n78), .Z(\ML_int[1][15] ) );
  MUX2_X1 M1_0_14 ( .A(A[14]), .B(A[13]), .S(n77), .Z(\ML_int[1][14] ) );
  MUX2_X1 M1_0_13 ( .A(A[13]), .B(A[12]), .S(SH[0]), .Z(\ML_int[1][13] ) );
  MUX2_X1 M1_0_12 ( .A(A[12]), .B(A[11]), .S(SH[0]), .Z(\ML_int[1][12] ) );
  MUX2_X1 M1_0_11 ( .A(A[11]), .B(A[10]), .S(n78), .Z(\ML_int[1][11] ) );
  MUX2_X1 M1_0_10 ( .A(A[10]), .B(A[9]), .S(n78), .Z(\ML_int[1][10] ) );
  MUX2_X1 M1_0_9 ( .A(A[9]), .B(A[8]), .S(n77), .Z(\ML_int[1][9] ) );
  MUX2_X1 M1_0_8 ( .A(A[8]), .B(A[7]), .S(n77), .Z(\ML_int[1][8] ) );
  MUX2_X1 M1_0_7 ( .A(A[7]), .B(A[6]), .S(n77), .Z(\ML_int[1][7] ) );
  MUX2_X1 M1_0_6 ( .A(A[6]), .B(A[5]), .S(n77), .Z(\ML_int[1][6] ) );
  MUX2_X1 M1_0_5 ( .A(A[5]), .B(A[4]), .S(n77), .Z(\ML_int[1][5] ) );
  MUX2_X1 M1_0_4 ( .A(A[4]), .B(A[3]), .S(n77), .Z(\ML_int[1][4] ) );
  MUX2_X1 M1_0_3 ( .A(A[3]), .B(A[2]), .S(n77), .Z(\ML_int[1][3] ) );
  MUX2_X1 M1_0_2 ( .A(A[2]), .B(A[1]), .S(n77), .Z(\ML_int[1][2] ) );
  MUX2_X1 M1_0_1 ( .A(A[1]), .B(A[0]), .S(n77), .Z(\ML_int[1][1] ) );
  NOR2_X1 U3 ( .A1(n86), .A2(n8), .ZN(B[2]) );
  NOR2_X1 U4 ( .A1(n86), .A2(n7), .ZN(B[3]) );
  NOR2_X1 U5 ( .A1(n86), .A2(n6), .ZN(B[4]) );
  NOR2_X1 U6 ( .A1(n86), .A2(n5), .ZN(B[5]) );
  NOR2_X1 U7 ( .A1(n86), .A2(n4), .ZN(B[6]) );
  NOR2_X1 U8 ( .A1(n86), .A2(n3), .ZN(B[7]) );
  INV_X1 U9 ( .A(n8), .ZN(\ML_int[4][2] ) );
  INV_X1 U10 ( .A(n6), .ZN(\ML_int[4][4] ) );
  INV_X1 U11 ( .A(n5), .ZN(\ML_int[4][5] ) );
  INV_X1 U12 ( .A(n4), .ZN(\ML_int[4][6] ) );
  INV_X1 U13 ( .A(n10), .ZN(\ML_int[4][0] ) );
  INV_X1 U14 ( .A(n9), .ZN(\ML_int[4][1] ) );
  INV_X1 U15 ( .A(n7), .ZN(\ML_int[4][3] ) );
  INV_X1 U16 ( .A(n3), .ZN(\ML_int[4][7] ) );
  NOR2_X1 U17 ( .A1(n86), .A2(n10), .ZN(B[0]) );
  NOR2_X1 U18 ( .A1(n86), .A2(n9), .ZN(B[1]) );
  INV_X1 U19 ( .A(n85), .ZN(n83) );
  INV_X1 U20 ( .A(n85), .ZN(n84) );
  NAND2_X1 U21 ( .A1(\ML_int[3][0] ), .A2(n85), .ZN(n10) );
  NAND2_X1 U22 ( .A1(\ML_int[3][1] ), .A2(n85), .ZN(n9) );
  NAND2_X1 U23 ( .A1(\ML_int[3][2] ), .A2(n85), .ZN(n8) );
  NAND2_X1 U24 ( .A1(\ML_int[3][3] ), .A2(n85), .ZN(n7) );
  NAND2_X1 U25 ( .A1(\ML_int[3][4] ), .A2(n85), .ZN(n6) );
  NAND2_X1 U26 ( .A1(\ML_int[3][5] ), .A2(n85), .ZN(n5) );
  NAND2_X1 U27 ( .A1(\ML_int[3][6] ), .A2(n85), .ZN(n4) );
  NAND2_X1 U28 ( .A1(\ML_int[3][7] ), .A2(n85), .ZN(n3) );
  AND2_X1 U29 ( .A1(\ML_int[4][8] ), .A2(n87), .ZN(B[8]) );
  AND2_X1 U30 ( .A1(\ML_int[4][9] ), .A2(n87), .ZN(B[9]) );
  AND2_X1 U31 ( .A1(\ML_int[4][10] ), .A2(n87), .ZN(B[10]) );
  AND2_X1 U32 ( .A1(\ML_int[4][11] ), .A2(n87), .ZN(B[11]) );
  AND2_X1 U33 ( .A1(\ML_int[4][12] ), .A2(n87), .ZN(B[12]) );
  AND2_X1 U34 ( .A1(\ML_int[4][13] ), .A2(n87), .ZN(B[13]) );
  AND2_X1 U35 ( .A1(\ML_int[4][14] ), .A2(n87), .ZN(B[14]) );
  AND2_X1 U36 ( .A1(\ML_int[4][15] ), .A2(n87), .ZN(B[15]) );
  INV_X1 U37 ( .A(n79), .ZN(n77) );
  INV_X1 U38 ( .A(n79), .ZN(n78) );
  INV_X1 U39 ( .A(n82), .ZN(n81) );
  INV_X1 U40 ( .A(SH[4]), .ZN(n87) );
  AND2_X1 U41 ( .A1(\ML_int[2][0] ), .A2(n82), .ZN(\ML_int[3][0] ) );
  AND2_X1 U42 ( .A1(\ML_int[2][1] ), .A2(n82), .ZN(\ML_int[3][1] ) );
  AND2_X1 U43 ( .A1(\ML_int[2][2] ), .A2(n82), .ZN(\ML_int[3][2] ) );
  AND2_X1 U44 ( .A1(\ML_int[2][3] ), .A2(n82), .ZN(\ML_int[3][3] ) );
  AND2_X1 U45 ( .A1(\ML_int[1][0] ), .A2(n76), .ZN(\ML_int[2][0] ) );
  AND2_X1 U46 ( .A1(\ML_int[1][1] ), .A2(n76), .ZN(\ML_int[2][1] ) );
  INV_X1 U47 ( .A(SH[2]), .ZN(n82) );
  INV_X1 U48 ( .A(SH[0]), .ZN(n79) );
  INV_X1 U49 ( .A(SH[1]), .ZN(n76) );
  INV_X1 U50 ( .A(n76), .ZN(n74) );
  INV_X1 U51 ( .A(n76), .ZN(n75) );
  AND2_X1 U52 ( .A1(A[0]), .A2(n79), .ZN(\ML_int[1][0] ) );
  INV_X1 U53 ( .A(n82), .ZN(n80) );
  INV_X1 U54 ( .A(SH[3]), .ZN(n85) );
  INV_X1 U55 ( .A(n87), .ZN(n86) );
endmodule


module FA_65 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3, n15, n16;

  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n2), .ZN(n16) );
  INV_X1 U2 ( .A(n3), .ZN(Co) );
  CLKBUF_X1 U3 ( .A(Ci), .Z(n15) );
  AOI22_X1 U5 ( .A1(B), .A2(A), .B1(n2), .B2(n15), .ZN(n3) );
  XNOR2_X1 U6 ( .A(Ci), .B(n16), .ZN(S) );
endmodule


module FA_66 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n26, n27, n29, n30, n31, n32, n33;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(n29) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n31) );
  NOR2_X1 U3 ( .A1(n29), .A2(n30), .ZN(n26) );
  AOI21_X1 U4 ( .B1(n32), .B2(Ci), .A(n26), .ZN(n27) );
  INV_X1 U5 ( .A(n27), .ZN(Co) );
  NAND2_X1 U6 ( .A1(n31), .A2(n29), .ZN(n32) );
  INV_X1 U7 ( .A(n32), .ZN(n30) );
  XNOR2_X1 U8 ( .A(n33), .B(n31), .ZN(S) );
  CLKBUF_X1 U9 ( .A(Ci), .Z(n33) );
endmodule


module FA_67 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net195774, net195771, n25, n26, n27, n28, n29, n30;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(n25) );
  NOR2_X1 U2 ( .A1(n28), .A2(n29), .ZN(n27) );
  INV_X1 U3 ( .A(n30), .ZN(n29) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n30) );
  XNOR2_X1 U5 ( .A(net195771), .B(n30), .ZN(S) );
  INV_X1 U6 ( .A(n25), .ZN(n28) );
  AOI21_X1 U7 ( .B1(n26), .B2(n25), .A(n27), .ZN(Co) );
  INV_X1 U8 ( .A(Ci), .ZN(n26) );
  CLKBUF_X1 U9 ( .A(n26), .Z(net195774) );
  INV_X1 U10 ( .A(net195774), .ZN(net195771) );
endmodule


module FA_68 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103612, n27, n28, n29, n30, n31, n32, n33, n34;
  assign Co = net103612;

  NOR2_X1 U1 ( .A1(n30), .A2(n31), .ZN(n29) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n27) );
  INV_X1 U3 ( .A(n32), .ZN(n31) );
  XNOR2_X1 U4 ( .A(B), .B(A), .ZN(n32) );
  XNOR2_X1 U5 ( .A(n33), .B(n32), .ZN(S) );
  INV_X1 U6 ( .A(n27), .ZN(n30) );
  INV_X1 U7 ( .A(Ci), .ZN(n28) );
  INV_X1 U8 ( .A(n34), .ZN(n33) );
  AOI21_X1 U9 ( .B1(n28), .B2(n27), .A(n29), .ZN(net103612) );
  CLKBUF_X1 U10 ( .A(n28), .Z(n34) );
endmodule


module FA_69 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103615, n30, n31, n32, n33, n34, n35, n36, n37;
  assign Co = net103615;

  NOR2_X1 U1 ( .A1(n35), .A2(n36), .ZN(n34) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n32) );
  INV_X1 U3 ( .A(n37), .ZN(n36) );
  XNOR2_X1 U4 ( .A(A), .B(B), .ZN(n37) );
  XNOR2_X1 U5 ( .A(n31), .B(n37), .ZN(S) );
  CLKBUF_X1 U6 ( .A(n33), .Z(n30) );
  INV_X1 U7 ( .A(n30), .ZN(n31) );
  INV_X1 U8 ( .A(n32), .ZN(n35) );
  AOI21_X1 U9 ( .B1(n33), .B2(n32), .A(n34), .ZN(net103615) );
  INV_X1 U10 ( .A(Ci), .ZN(n33) );
endmodule


module FA_70 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103618, net198326, net198323, n25, n26, n27, n28;
  assign Co = net103618;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(n26) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n28) );
  XNOR2_X1 U3 ( .A(net198323), .B(n28), .ZN(S) );
  AND2_X1 U4 ( .A1(n28), .A2(n26), .ZN(n25) );
  AOI21_X1 U5 ( .B1(n27), .B2(n26), .A(n25), .ZN(net103618) );
  INV_X1 U6 ( .A(Ci), .ZN(n27) );
  CLKBUF_X1 U7 ( .A(n27), .Z(net198326) );
  INV_X1 U8 ( .A(net198326), .ZN(net198323) );
endmodule


module FA_71 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103621, net196874, net196871, n24, n25, n26, n27;
  assign Co = net103621;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(n25) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n27) );
  XNOR2_X1 U3 ( .A(net196871), .B(n27), .ZN(S) );
  AND2_X1 U4 ( .A1(n27), .A2(n25), .ZN(n24) );
  AOI21_X1 U5 ( .B1(n26), .B2(n25), .A(n24), .ZN(net103621) );
  INV_X1 U6 ( .A(Ci), .ZN(n26) );
  CLKBUF_X1 U7 ( .A(n26), .Z(net196874) );
  INV_X1 U8 ( .A(net196874), .ZN(net196871) );
endmodule


module FA_72 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103624, net196650, net196647, n26, n27, n28, n29;
  assign Co = net103624;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(n27) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n29) );
  XNOR2_X1 U3 ( .A(net196647), .B(n29), .ZN(S) );
  AND2_X1 U4 ( .A1(n29), .A2(n27), .ZN(n26) );
  AOI21_X1 U5 ( .B1(n28), .B2(n27), .A(n26), .ZN(net103624) );
  INV_X1 U6 ( .A(Ci), .ZN(n28) );
  CLKBUF_X1 U7 ( .A(n28), .Z(net196650) );
  INV_X1 U8 ( .A(net196650), .ZN(net196647) );
endmodule


module FA_73 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103627, n30, n31, n32, n33, n34, n35;
  assign Co = net103627;

  XNOR2_X1 U1 ( .A(n32), .B(n35), .ZN(S) );
  AND2_X1 U2 ( .A1(n35), .A2(n33), .ZN(n30) );
  XNOR2_X1 U3 ( .A(A), .B(B), .ZN(n35) );
  NAND2_X1 U4 ( .A1(A), .A2(B), .ZN(n33) );
  AOI21_X1 U5 ( .B1(n34), .B2(n33), .A(n30), .ZN(net103627) );
  CLKBUF_X1 U6 ( .A(n34), .Z(n31) );
  INV_X1 U7 ( .A(n31), .ZN(n32) );
  INV_X1 U8 ( .A(Ci), .ZN(n34) );
endmodule


module FA_74 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103630, net197100, net197097, n25, n26, n27, n28, n29, n30;
  assign Co = net103630;

  NOR2_X1 U1 ( .A1(n28), .A2(n29), .ZN(n27) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n30) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n25) );
  INV_X1 U4 ( .A(n30), .ZN(n29) );
  XNOR2_X1 U5 ( .A(net197097), .B(n30), .ZN(S) );
  INV_X1 U6 ( .A(n25), .ZN(n28) );
  AOI21_X1 U7 ( .B1(n26), .B2(n25), .A(n27), .ZN(net103630) );
  INV_X1 U8 ( .A(Ci), .ZN(n26) );
  CLKBUF_X1 U9 ( .A(n26), .Z(net197100) );
  INV_X1 U10 ( .A(net197100), .ZN(net197097) );
endmodule


module FA_75 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103633, n32, n33, n34, n35, n36, n37;
  assign Co = net103633;

  XNOR2_X1 U1 ( .A(n34), .B(n37), .ZN(S) );
  AND2_X1 U2 ( .A1(n37), .A2(n35), .ZN(n32) );
  CLKBUF_X1 U3 ( .A(n36), .Z(n33) );
  INV_X1 U4 ( .A(n33), .ZN(n34) );
  XNOR2_X1 U5 ( .A(A), .B(B), .ZN(n37) );
  NAND2_X1 U6 ( .A1(A), .A2(B), .ZN(n35) );
  AOI21_X1 U7 ( .B1(n36), .B2(n35), .A(n32), .ZN(net103633) );
  INV_X1 U8 ( .A(Ci), .ZN(n36) );
endmodule


module FA_76 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103636, net197536, net197533, n25, n26, n27, n28, n29, n30;
  assign Co = net103636;

  NOR2_X1 U1 ( .A1(n28), .A2(n29), .ZN(n27) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n30) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n25) );
  INV_X1 U4 ( .A(n30), .ZN(n29) );
  XNOR2_X1 U5 ( .A(net197533), .B(n30), .ZN(S) );
  INV_X1 U6 ( .A(n25), .ZN(n28) );
  AOI21_X1 U7 ( .B1(n26), .B2(n25), .A(n27), .ZN(net103636) );
  INV_X1 U8 ( .A(Ci), .ZN(n26) );
  CLKBUF_X1 U9 ( .A(n26), .Z(net197536) );
  INV_X1 U10 ( .A(net197536), .ZN(net197533) );
endmodule


module FA_77 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n26, n27, n28, n29, n30, n31, n32, n33;

  NOR2_X1 U1 ( .A1(n31), .A2(n32), .ZN(n30) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n33) );
  NAND2_X1 U3 ( .A1(A), .A2(B), .ZN(n28) );
  INV_X1 U4 ( .A(n33), .ZN(n32) );
  XNOR2_X1 U5 ( .A(n27), .B(n33), .ZN(S) );
  CLKBUF_X1 U6 ( .A(n29), .Z(n26) );
  INV_X1 U7 ( .A(n26), .ZN(n27) );
  INV_X1 U8 ( .A(n28), .ZN(n31) );
  AOI21_X1 U9 ( .B1(n29), .B2(n28), .A(n30), .ZN(Co) );
  INV_X1 U10 ( .A(Ci), .ZN(n29) );
endmodule


module FA_78 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n26, n27, n29;

  XOR2_X1 U3 ( .A(n29), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(n26) );
  AOI21_X1 U2 ( .B1(Ci), .B2(n2), .A(n26), .ZN(n27) );
  INV_X1 U5 ( .A(n27), .ZN(Co) );
  CLKBUF_X1 U6 ( .A(Ci), .Z(n29) );
endmodule


module FA_79 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n27, n28, n30, n31, n32, n33, n34, n35, n36;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(n31) );
  XNOR2_X1 U2 ( .A(A), .B(B), .ZN(n35) );
  INV_X1 U3 ( .A(n35), .ZN(n34) );
  XNOR2_X1 U4 ( .A(n36), .B(n35), .ZN(S) );
  NOR2_X1 U5 ( .A1(n31), .A2(n32), .ZN(n27) );
  AOI21_X1 U6 ( .B1(Ci), .B2(n30), .A(n27), .ZN(n28) );
  INV_X1 U7 ( .A(n28), .ZN(Co) );
  INV_X1 U8 ( .A(n32), .ZN(n30) );
  NOR2_X1 U9 ( .A1(n33), .A2(n34), .ZN(n32) );
  INV_X1 U10 ( .A(n31), .ZN(n33) );
  CLKBUF_X1 U11 ( .A(Ci), .Z(n36) );
endmodule


module FA_80 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n25, n26, n28, n29, n30, n31, n32;

  XNOR2_X1 U1 ( .A(A), .B(B), .ZN(n30) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n28) );
  XNOR2_X1 U3 ( .A(n32), .B(n30), .ZN(S) );
  NAND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(Co) );
  OR2_X1 U5 ( .A1(n28), .A2(n29), .ZN(n25) );
  NAND2_X1 U6 ( .A1(Ci), .A2(n31), .ZN(n26) );
  NAND2_X1 U7 ( .A1(n30), .A2(n28), .ZN(n31) );
  INV_X1 U8 ( .A(n31), .ZN(n29) );
  CLKBUF_X1 U9 ( .A(Ci), .Z(n32) );
endmodule


module FA_81 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103651, n27, n28, n29, n30, n31, n32;
  assign Co = net103651;

  XNOR2_X1 U1 ( .A(B), .B(A), .ZN(n30) );
  NAND2_X1 U2 ( .A1(A), .A2(B), .ZN(n28) );
  XNOR2_X1 U3 ( .A(n31), .B(n30), .ZN(S) );
  AND2_X1 U4 ( .A1(n30), .A2(n28), .ZN(n27) );
  AOI21_X1 U5 ( .B1(n29), .B2(n28), .A(n27), .ZN(net103651) );
  INV_X1 U6 ( .A(Ci), .ZN(n29) );
  INV_X1 U7 ( .A(n32), .ZN(n31) );
  CLKBUF_X1 U8 ( .A(n29), .Z(n32) );
endmodule


module FA_82 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net195854, net195851, n25, n26, n27, n28;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(n26) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n28) );
  XNOR2_X1 U3 ( .A(net195851), .B(n28), .ZN(S) );
  AND2_X1 U4 ( .A1(n28), .A2(n26), .ZN(n25) );
  AOI21_X1 U5 ( .B1(n27), .B2(n26), .A(n25), .ZN(Co) );
  INV_X1 U6 ( .A(Ci), .ZN(n27) );
  CLKBUF_X1 U7 ( .A(n27), .Z(net195854) );
  INV_X1 U8 ( .A(net195854), .ZN(net195851) );
endmodule


module FA_83 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103657, n24, n25, n26, n27, n28, n29;
  assign Co = net103657;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(n25) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n27) );
  XNOR2_X1 U3 ( .A(n28), .B(n27), .ZN(S) );
  AND2_X1 U4 ( .A1(n27), .A2(n25), .ZN(n24) );
  AOI21_X1 U5 ( .B1(n26), .B2(n25), .A(n24), .ZN(net103657) );
  INV_X1 U6 ( .A(Ci), .ZN(n26) );
  INV_X1 U7 ( .A(n29), .ZN(n28) );
  CLKBUF_X1 U8 ( .A(n26), .Z(n29) );
endmodule


module FA_84 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   net103660, n29, n30, n31, n32, n33, n34;
  assign Co = net103660;

  NAND2_X1 U1 ( .A1(A), .A2(B), .ZN(n31) );
  XNOR2_X1 U2 ( .A(B), .B(A), .ZN(n33) );
  XNOR2_X1 U3 ( .A(n34), .B(n33), .ZN(S) );
  CLKBUF_X1 U4 ( .A(n32), .Z(n29) );
  AND2_X1 U5 ( .A1(n33), .A2(n31), .ZN(n30) );
  AOI21_X1 U6 ( .B1(n32), .B2(n31), .A(n30), .ZN(net103660) );
  INV_X1 U7 ( .A(Ci), .ZN(n32) );
  INV_X1 U8 ( .A(n29), .ZN(n34) );
endmodule


module FA_85 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n3, n28, n29, n31;

  XOR2_X1 U3 ( .A(n31), .B(n3), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n3) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(n28) );
  AOI21_X1 U2 ( .B1(Ci), .B2(n3), .A(n28), .ZN(n29) );
  INV_X1 U5 ( .A(n29), .ZN(Co) );
  CLKBUF_X1 U6 ( .A(Ci), .Z(n31) );
endmodule


module FA_86 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n25, n26, n28;

  XOR2_X1 U3 ( .A(n28), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(n25) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n2), .ZN(n26) );
  NAND2_X1 U5 ( .A1(n26), .A2(n25), .ZN(Co) );
  CLKBUF_X1 U6 ( .A(Ci), .Z(n28) );
endmodule


module FA_87 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n24, n25, n27;

  XOR2_X1 U3 ( .A(n27), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(n24) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n2), .ZN(n25) );
  NAND2_X1 U5 ( .A1(n25), .A2(n24), .ZN(Co) );
  CLKBUF_X1 U6 ( .A(Ci), .Z(n27) );
endmodule


module FA_88 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n24, n25, n27;

  XOR2_X1 U3 ( .A(n27), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(n24) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n2), .ZN(n25) );
  NAND2_X1 U5 ( .A1(n25), .A2(n24), .ZN(Co) );
  CLKBUF_X1 U6 ( .A(Ci), .Z(n27) );
endmodule


module FA_89 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n22, n23, n25;

  XOR2_X1 U3 ( .A(n25), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(n22) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n2), .ZN(n23) );
  NAND2_X1 U5 ( .A1(n23), .A2(n22), .ZN(Co) );
  CLKBUF_X1 U6 ( .A(Ci), .Z(n25) );
endmodule


module FA_90 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n21, n22, n24;

  XOR2_X1 U3 ( .A(n24), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(n21) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n2), .ZN(n22) );
  NAND2_X1 U5 ( .A1(n22), .A2(n21), .ZN(Co) );
  CLKBUF_X1 U6 ( .A(Ci), .Z(n24) );
endmodule


module FA_91 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n22, n23, n24, n26;

  XOR2_X1 U3 ( .A(n26), .B(n2), .Z(S) );
  INV_X1 U1 ( .A(B), .ZN(n22) );
  XNOR2_X1 U2 ( .A(A), .B(n22), .ZN(n2) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n23) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n2), .ZN(n24) );
  NAND2_X1 U6 ( .A1(n23), .A2(n24), .ZN(Co) );
  CLKBUF_X1 U7 ( .A(Ci), .Z(n26) );
endmodule


module FA_92 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n22, n23, n24, n26;

  XOR2_X1 U3 ( .A(n26), .B(n2), .Z(S) );
  INV_X1 U1 ( .A(B), .ZN(n22) );
  XNOR2_X1 U2 ( .A(A), .B(n22), .ZN(n2) );
  NAND2_X1 U4 ( .A1(B), .A2(A), .ZN(n23) );
  NAND2_X1 U5 ( .A1(Ci), .A2(n2), .ZN(n24) );
  NAND2_X1 U6 ( .A1(n24), .A2(n23), .ZN(Co) );
  CLKBUF_X1 U7 ( .A(Ci), .Z(n26) );
endmodule


module FA_93 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n25, n26, n28, n29;

  XOR2_X1 U3 ( .A(n29), .B(n2), .Z(S) );
  INV_X1 U1 ( .A(B), .ZN(n28) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n25) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n2), .ZN(n26) );
  NAND2_X1 U5 ( .A1(n25), .A2(n26), .ZN(Co) );
  XNOR2_X1 U6 ( .A(A), .B(n28), .ZN(n2) );
  CLKBUF_X1 U7 ( .A(Ci), .Z(n29) );
endmodule


module FA_94 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n26, n27, n29, n30;

  XOR2_X1 U3 ( .A(n30), .B(n2), .Z(S) );
  INV_X1 U1 ( .A(B), .ZN(n29) );
  NAND2_X1 U2 ( .A1(B), .A2(A), .ZN(n26) );
  NAND2_X1 U4 ( .A1(Ci), .A2(n2), .ZN(n27) );
  NAND2_X1 U5 ( .A1(n26), .A2(n27), .ZN(Co) );
  XNOR2_X1 U6 ( .A(A), .B(n29), .ZN(n2) );
  CLKBUF_X1 U7 ( .A(Ci), .Z(n30) );
endmodule


module FA_95 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n31, n32, n34, n35;

  XOR2_X1 U3 ( .A(n35), .B(n2), .Z(S) );
  NAND2_X1 U1 ( .A1(B), .A2(A), .ZN(n31) );
  NAND2_X1 U2 ( .A1(Ci), .A2(n2), .ZN(n32) );
  NAND2_X1 U4 ( .A1(n31), .A2(n32), .ZN(Co) );
  INV_X1 U5 ( .A(B), .ZN(n34) );
  XNOR2_X1 U6 ( .A(A), .B(n34), .ZN(n2) );
  CLKBUF_X1 U7 ( .A(Ci), .Z(n35) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n28, n29, n31, n32, n33;

  XOR2_X1 U3 ( .A(Ci), .B(n33), .Z(S) );
  NAND2_X1 U1 ( .A1(B), .A2(n32), .ZN(n28) );
  NAND2_X1 U2 ( .A1(n2), .A2(Ci), .ZN(n29) );
  NAND2_X1 U4 ( .A1(n28), .A2(n29), .ZN(Co) );
  INV_X1 U5 ( .A(B), .ZN(n31) );
  XNOR2_X1 U6 ( .A(A), .B(n31), .ZN(n2) );
  CLKBUF_X1 U7 ( .A(A), .Z(n32) );
  CLKBUF_X1 U8 ( .A(n2), .Z(n33) );
endmodule


module MUX_6to1_n32 ( A, B, C, D, E, F, S, Y );
  input [31:0] A;
  input [31:0] B;
  input [31:0] C;
  input [31:0] D;
  input [31:0] E;
  input [31:0] F;
  input [2:0] S;
  output [31:0] Y;
  wire   n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194;

  BUF_X1 U1 ( .A(n188), .Z(n189) );
  BUF_X1 U2 ( .A(n188), .Z(n190) );
  BUF_X1 U3 ( .A(n188), .Z(n191) );
  BUF_X1 U4 ( .A(n11), .Z(n176) );
  BUF_X1 U5 ( .A(n8), .Z(n186) );
  BUF_X1 U6 ( .A(n11), .Z(n177) );
  BUF_X1 U7 ( .A(n8), .Z(n185) );
  BUF_X1 U8 ( .A(n11), .Z(n178) );
  BUF_X1 U9 ( .A(n8), .Z(n187) );
  BUF_X1 U10 ( .A(n7), .Z(n188) );
  NOR4_X1 U11 ( .A1(n176), .A2(n182), .A3(n179), .A4(n74), .ZN(n7) );
  OR2_X1 U12 ( .A1(n194), .A2(n187), .ZN(n74) );
  BUF_X1 U13 ( .A(n10), .Z(n179) );
  BUF_X1 U14 ( .A(n10), .Z(n180) );
  BUF_X1 U15 ( .A(n9), .Z(n182) );
  BUF_X1 U16 ( .A(n9), .Z(n183) );
  BUF_X1 U17 ( .A(n6), .Z(n193) );
  BUF_X1 U18 ( .A(n6), .Z(n192) );
  NOR3_X1 U19 ( .A1(n77), .A2(S[2]), .A3(n75), .ZN(n11) );
  NOR3_X1 U20 ( .A1(S[0]), .A2(S[2]), .A3(n75), .ZN(n8) );
  BUF_X1 U21 ( .A(n6), .Z(n194) );
  BUF_X1 U22 ( .A(n10), .Z(n181) );
  BUF_X1 U23 ( .A(n9), .Z(n184) );
  INV_X1 U24 ( .A(S[0]), .ZN(n77) );
  INV_X1 U25 ( .A(S[2]), .ZN(n76) );
  AOI222_X1 U26 ( .A1(E[2]), .A2(n182), .B1(B[2]), .B2(n179), .C1(D[2]), .C2(
        n176), .ZN(n28) );
  AOI222_X1 U27 ( .A1(E[5]), .A2(n182), .B1(B[5]), .B2(n179), .C1(D[5]), .C2(
        n176), .ZN(n18) );
  AOI222_X1 U28 ( .A1(E[30]), .A2(n182), .B1(B[30]), .B2(n179), .C1(D[30]), 
        .C2(n176), .ZN(n26) );
  AOI222_X1 U29 ( .A1(E[6]), .A2(n182), .B1(B[6]), .B2(n179), .C1(D[6]), .C2(
        n176), .ZN(n16) );
  AOI222_X1 U30 ( .A1(E[7]), .A2(n182), .B1(B[7]), .B2(n179), .C1(D[7]), .C2(
        n176), .ZN(n14) );
  AOI222_X1 U31 ( .A1(E[4]), .A2(n182), .B1(B[4]), .B2(n179), .C1(D[4]), .C2(
        n176), .ZN(n20) );
  AOI222_X1 U32 ( .A1(E[31]), .A2(n182), .B1(B[31]), .B2(n179), .C1(D[31]), 
        .C2(n176), .ZN(n24) );
  AOI222_X1 U33 ( .A1(E[3]), .A2(n182), .B1(B[3]), .B2(n179), .C1(D[3]), .C2(
        n176), .ZN(n22) );
  AOI222_X1 U34 ( .A1(E[23]), .A2(n183), .B1(B[23]), .B2(n180), .C1(D[23]), 
        .C2(n177), .ZN(n42) );
  AOI222_X1 U35 ( .A1(E[1]), .A2(n183), .B1(B[1]), .B2(n180), .C1(D[1]), .C2(
        n177), .ZN(n50) );
  AOI222_X1 U36 ( .A1(E[24]), .A2(n183), .B1(B[24]), .B2(n180), .C1(D[24]), 
        .C2(n177), .ZN(n40) );
  AOI222_X1 U37 ( .A1(E[25]), .A2(n183), .B1(B[25]), .B2(n180), .C1(D[25]), 
        .C2(n177), .ZN(n38) );
  AOI222_X1 U38 ( .A1(E[27]), .A2(n183), .B1(B[27]), .B2(n180), .C1(D[27]), 
        .C2(n177), .ZN(n34) );
  AOI222_X1 U39 ( .A1(E[28]), .A2(n183), .B1(B[28]), .B2(n180), .C1(D[28]), 
        .C2(n177), .ZN(n32) );
  AOI222_X1 U40 ( .A1(E[0]), .A2(n182), .B1(B[0]), .B2(n179), .C1(D[0]), .C2(
        n176), .ZN(n72) );
  AOI222_X1 U41 ( .A1(E[19]), .A2(n183), .B1(B[19]), .B2(n180), .C1(D[19]), 
        .C2(n177), .ZN(n52) );
  AOI222_X1 U42 ( .A1(E[26]), .A2(n183), .B1(B[26]), .B2(n180), .C1(D[26]), 
        .C2(n177), .ZN(n36) );
  AOI222_X1 U43 ( .A1(E[8]), .A2(n182), .B1(B[8]), .B2(n179), .C1(D[8]), .C2(
        n176), .ZN(n12) );
  AOI222_X1 U44 ( .A1(E[9]), .A2(n183), .B1(B[9]), .B2(n180), .C1(D[9]), .C2(
        n177), .ZN(n4) );
  AOI222_X1 U45 ( .A1(E[29]), .A2(n182), .B1(B[29]), .B2(n179), .C1(D[29]), 
        .C2(n176), .ZN(n30) );
  AOI222_X1 U46 ( .A1(E[20]), .A2(n183), .B1(B[20]), .B2(n180), .C1(D[20]), 
        .C2(n177), .ZN(n48) );
  AOI222_X1 U47 ( .A1(E[21]), .A2(n183), .B1(B[21]), .B2(n180), .C1(D[21]), 
        .C2(n177), .ZN(n46) );
  AOI222_X1 U48 ( .A1(E[22]), .A2(n183), .B1(B[22]), .B2(n180), .C1(D[22]), 
        .C2(n177), .ZN(n44) );
  AOI222_X1 U49 ( .A1(E[10]), .A2(n184), .B1(B[10]), .B2(n181), .C1(D[10]), 
        .C2(n178), .ZN(n70) );
  AOI222_X1 U50 ( .A1(E[11]), .A2(n184), .B1(B[11]), .B2(n181), .C1(D[11]), 
        .C2(n178), .ZN(n68) );
  AOI222_X1 U51 ( .A1(E[12]), .A2(n184), .B1(B[12]), .B2(n181), .C1(D[12]), 
        .C2(n178), .ZN(n66) );
  AOI222_X1 U52 ( .A1(E[13]), .A2(n184), .B1(B[13]), .B2(n181), .C1(D[13]), 
        .C2(n178), .ZN(n64) );
  AOI222_X1 U53 ( .A1(E[14]), .A2(n184), .B1(B[14]), .B2(n181), .C1(D[14]), 
        .C2(n178), .ZN(n62) );
  AOI222_X1 U54 ( .A1(E[15]), .A2(n184), .B1(B[15]), .B2(n181), .C1(D[15]), 
        .C2(n178), .ZN(n60) );
  AOI222_X1 U55 ( .A1(E[16]), .A2(n184), .B1(B[16]), .B2(n181), .C1(D[16]), 
        .C2(n178), .ZN(n58) );
  AOI222_X1 U56 ( .A1(E[17]), .A2(n184), .B1(B[17]), .B2(n181), .C1(D[17]), 
        .C2(n178), .ZN(n56) );
  AOI222_X1 U57 ( .A1(E[18]), .A2(n184), .B1(B[18]), .B2(n181), .C1(D[18]), 
        .C2(n178), .ZN(n54) );
  NOR3_X1 U58 ( .A1(S[1]), .A2(S[2]), .A3(n77), .ZN(n10) );
  NOR3_X1 U59 ( .A1(S[0]), .A2(S[1]), .A3(n76), .ZN(n9) );
  NOR3_X1 U60 ( .A1(n76), .A2(S[1]), .A3(n77), .ZN(n6) );
  INV_X1 U61 ( .A(S[1]), .ZN(n75) );
  NAND2_X1 U62 ( .A1(n50), .A2(n51), .ZN(Y[1]) );
  AOI222_X1 U63 ( .A1(F[1]), .A2(n193), .B1(A[1]), .B2(n189), .C1(C[1]), .C2(
        n186), .ZN(n51) );
  NAND2_X1 U64 ( .A1(n40), .A2(n41), .ZN(Y[24]) );
  AOI222_X1 U65 ( .A1(F[24]), .A2(n193), .B1(A[24]), .B2(n190), .C1(C[24]), 
        .C2(n186), .ZN(n41) );
  NAND2_X1 U66 ( .A1(n38), .A2(n39), .ZN(Y[25]) );
  AOI222_X1 U67 ( .A1(F[25]), .A2(n193), .B1(A[25]), .B2(n190), .C1(C[25]), 
        .C2(n186), .ZN(n39) );
  NAND2_X1 U68 ( .A1(n34), .A2(n35), .ZN(Y[27]) );
  AOI222_X1 U69 ( .A1(F[27]), .A2(n193), .B1(A[27]), .B2(n190), .C1(C[27]), 
        .C2(n186), .ZN(n35) );
  NAND2_X1 U70 ( .A1(n32), .A2(n33), .ZN(Y[28]) );
  AOI222_X1 U71 ( .A1(F[28]), .A2(n193), .B1(A[28]), .B2(n190), .C1(C[28]), 
        .C2(n185), .ZN(n33) );
  NAND2_X1 U72 ( .A1(n28), .A2(n29), .ZN(Y[2]) );
  AOI222_X1 U73 ( .A1(F[2]), .A2(n192), .B1(A[2]), .B2(n190), .C1(C[2]), .C2(
        n185), .ZN(n29) );
  NAND2_X1 U74 ( .A1(n18), .A2(n19), .ZN(Y[5]) );
  AOI222_X1 U75 ( .A1(F[5]), .A2(n192), .B1(A[5]), .B2(n191), .C1(C[5]), .C2(
        n185), .ZN(n19) );
  NAND2_X1 U76 ( .A1(n26), .A2(n27), .ZN(Y[30]) );
  AOI222_X1 U77 ( .A1(F[30]), .A2(n192), .B1(A[30]), .B2(n190), .C1(C[30]), 
        .C2(n185), .ZN(n27) );
  NAND2_X1 U78 ( .A1(n16), .A2(n17), .ZN(Y[6]) );
  AOI222_X1 U79 ( .A1(F[6]), .A2(n192), .B1(A[6]), .B2(n191), .C1(C[6]), .C2(
        n185), .ZN(n17) );
  NAND2_X1 U80 ( .A1(n14), .A2(n15), .ZN(Y[7]) );
  AOI222_X1 U81 ( .A1(F[7]), .A2(n192), .B1(A[7]), .B2(n191), .C1(C[7]), .C2(
        n185), .ZN(n15) );
  NAND2_X1 U82 ( .A1(n20), .A2(n21), .ZN(Y[4]) );
  AOI222_X1 U83 ( .A1(F[4]), .A2(n192), .B1(A[4]), .B2(n191), .C1(C[4]), .C2(
        n185), .ZN(n21) );
  NAND2_X1 U84 ( .A1(n24), .A2(n25), .ZN(Y[31]) );
  AOI222_X1 U85 ( .A1(F[31]), .A2(n192), .B1(A[31]), .B2(n191), .C1(C[31]), 
        .C2(n185), .ZN(n25) );
  NAND2_X1 U86 ( .A1(n22), .A2(n23), .ZN(Y[3]) );
  AOI222_X1 U87 ( .A1(F[3]), .A2(n192), .B1(A[3]), .B2(n191), .C1(C[3]), .C2(
        n185), .ZN(n23) );
  NAND2_X1 U88 ( .A1(n42), .A2(n43), .ZN(Y[23]) );
  AOI222_X1 U89 ( .A1(F[23]), .A2(n193), .B1(A[23]), .B2(n190), .C1(C[23]), 
        .C2(n186), .ZN(n43) );
  NAND2_X1 U90 ( .A1(n72), .A2(n73), .ZN(Y[0]) );
  AOI222_X1 U91 ( .A1(F[0]), .A2(n194), .B1(A[0]), .B2(n189), .C1(C[0]), .C2(
        n187), .ZN(n73) );
  NAND2_X1 U92 ( .A1(n70), .A2(n71), .ZN(Y[10]) );
  AOI222_X1 U93 ( .A1(F[10]), .A2(n194), .B1(A[10]), .B2(n189), .C1(C[10]), 
        .C2(n187), .ZN(n71) );
  NAND2_X1 U94 ( .A1(n68), .A2(n69), .ZN(Y[11]) );
  AOI222_X1 U95 ( .A1(F[11]), .A2(n194), .B1(A[11]), .B2(n189), .C1(C[11]), 
        .C2(n187), .ZN(n69) );
  NAND2_X1 U96 ( .A1(n66), .A2(n67), .ZN(Y[12]) );
  AOI222_X1 U97 ( .A1(F[12]), .A2(n194), .B1(A[12]), .B2(n189), .C1(C[12]), 
        .C2(n187), .ZN(n67) );
  NAND2_X1 U98 ( .A1(n64), .A2(n65), .ZN(Y[13]) );
  AOI222_X1 U99 ( .A1(F[13]), .A2(n194), .B1(A[13]), .B2(n189), .C1(C[13]), 
        .C2(n187), .ZN(n65) );
  NAND2_X1 U100 ( .A1(n62), .A2(n63), .ZN(Y[14]) );
  AOI222_X1 U101 ( .A1(F[14]), .A2(n194), .B1(A[14]), .B2(n189), .C1(C[14]), 
        .C2(n187), .ZN(n63) );
  NAND2_X1 U102 ( .A1(n60), .A2(n61), .ZN(Y[15]) );
  AOI222_X1 U103 ( .A1(F[15]), .A2(n194), .B1(A[15]), .B2(n189), .C1(C[15]), 
        .C2(n187), .ZN(n61) );
  NAND2_X1 U104 ( .A1(n58), .A2(n59), .ZN(Y[16]) );
  AOI222_X1 U105 ( .A1(F[16]), .A2(n194), .B1(A[16]), .B2(n189), .C1(C[16]), 
        .C2(n187), .ZN(n59) );
  NAND2_X1 U106 ( .A1(n56), .A2(n57), .ZN(Y[17]) );
  AOI222_X1 U107 ( .A1(F[17]), .A2(n194), .B1(A[17]), .B2(n189), .C1(C[17]), 
        .C2(n186), .ZN(n57) );
  NAND2_X1 U108 ( .A1(n54), .A2(n55), .ZN(Y[18]) );
  AOI222_X1 U109 ( .A1(F[18]), .A2(n194), .B1(A[18]), .B2(n189), .C1(C[18]), 
        .C2(n186), .ZN(n55) );
  NAND2_X1 U110 ( .A1(n52), .A2(n53), .ZN(Y[19]) );
  AOI222_X1 U111 ( .A1(F[19]), .A2(n193), .B1(A[19]), .B2(n189), .C1(C[19]), 
        .C2(n186), .ZN(n53) );
  NAND2_X1 U112 ( .A1(n36), .A2(n37), .ZN(Y[26]) );
  AOI222_X1 U113 ( .A1(F[26]), .A2(n193), .B1(A[26]), .B2(n190), .C1(C[26]), 
        .C2(n186), .ZN(n37) );
  NAND2_X1 U114 ( .A1(n12), .A2(n13), .ZN(Y[8]) );
  AOI222_X1 U115 ( .A1(F[8]), .A2(n192), .B1(A[8]), .B2(n191), .C1(C[8]), .C2(
        n185), .ZN(n13) );
  NAND2_X1 U116 ( .A1(n4), .A2(n5), .ZN(Y[9]) );
  AOI222_X1 U117 ( .A1(F[9]), .A2(n192), .B1(A[9]), .B2(n191), .C1(C[9]), .C2(
        n185), .ZN(n5) );
  NAND2_X1 U118 ( .A1(n30), .A2(n31), .ZN(Y[29]) );
  AOI222_X1 U119 ( .A1(F[29]), .A2(n192), .B1(A[29]), .B2(n190), .C1(C[29]), 
        .C2(n185), .ZN(n31) );
  NAND2_X1 U120 ( .A1(n48), .A2(n49), .ZN(Y[20]) );
  AOI222_X1 U121 ( .A1(F[20]), .A2(n193), .B1(A[20]), .B2(n190), .C1(C[20]), 
        .C2(n186), .ZN(n49) );
  NAND2_X1 U122 ( .A1(n46), .A2(n47), .ZN(Y[21]) );
  AOI222_X1 U123 ( .A1(F[21]), .A2(n193), .B1(A[21]), .B2(n190), .C1(C[21]), 
        .C2(n186), .ZN(n47) );
  NAND2_X1 U124 ( .A1(n44), .A2(n45), .ZN(Y[22]) );
  AOI222_X1 U125 ( .A1(F[22]), .A2(n193), .B1(A[22]), .B2(n190), .C1(C[22]), 
        .C2(n186), .ZN(n45) );
endmodule


module MUX_2to1_n32 ( A, B, S, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input S;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108;
  assign Y[0] = N2;
  assign Y[1] = N3;
  assign Y[2] = N4;
  assign Y[3] = N5;
  assign Y[4] = N6;
  assign Y[5] = N7;
  assign Y[6] = N8;
  assign Y[7] = N9;
  assign Y[8] = N10;
  assign Y[9] = N11;
  assign Y[10] = N12;
  assign Y[11] = N13;
  assign Y[12] = N14;
  assign Y[13] = N15;
  assign Y[14] = N16;
  assign Y[15] = N17;
  assign Y[16] = N18;
  assign Y[17] = N19;
  assign Y[18] = N20;
  assign Y[19] = N21;
  assign Y[20] = N22;
  assign Y[21] = N23;
  assign Y[22] = N24;
  assign Y[23] = N25;
  assign Y[24] = N26;
  assign Y[25] = N27;
  assign Y[26] = N28;
  assign Y[27] = N29;
  assign Y[28] = N30;
  assign Y[29] = N31;
  assign Y[30] = N32;
  assign Y[31] = N33;

  BUF_X1 U1 ( .A(n97), .Z(n108) );
  BUF_X1 U2 ( .A(n97), .Z(n107) );
  INV_X1 U3 ( .A(n108), .ZN(n98) );
  BUF_X1 U4 ( .A(n96), .Z(n103) );
  BUF_X1 U5 ( .A(n95), .Z(n100) );
  CLKBUF_X1 U6 ( .A(n95), .Z(n101) );
  CLKBUF_X1 U7 ( .A(n95), .Z(n102) );
  CLKBUF_X1 U8 ( .A(n96), .Z(n105) );
  CLKBUF_X1 U9 ( .A(n96), .Z(n104) );
  BUF_X1 U10 ( .A(n97), .Z(n106) );
  BUF_X1 U11 ( .A(S), .Z(n97) );
  CLKBUF_X1 U12 ( .A(S), .Z(n96) );
  CLKBUF_X1 U13 ( .A(S), .Z(n95) );
  INV_X1 U14 ( .A(n40), .ZN(N4) );
  INV_X1 U15 ( .A(n37), .ZN(N7) );
  INV_X1 U16 ( .A(n42), .ZN(N32) );
  INV_X1 U17 ( .A(n36), .ZN(N8) );
  INV_X1 U18 ( .A(n34), .ZN(N9) );
  INV_X1 U19 ( .A(n38), .ZN(N6) );
  INV_X1 U20 ( .A(n41), .ZN(N33) );
  INV_X1 U21 ( .A(n39), .ZN(N5) );
  INV_X1 U22 ( .A(n50), .ZN(N25) );
  INV_X1 U23 ( .A(n45), .ZN(N3) );
  INV_X1 U24 ( .A(n49), .ZN(N26) );
  INV_X1 U25 ( .A(n48), .ZN(N27) );
  INV_X1 U26 ( .A(n46), .ZN(N29) );
  INV_X1 U27 ( .A(n44), .ZN(N30) );
  INV_X1 U28 ( .A(n56), .ZN(N2) );
  INV_X1 U29 ( .A(n54), .ZN(N21) );
  INV_X1 U30 ( .A(n47), .ZN(N28) );
  INV_X1 U31 ( .A(n66), .ZN(N10) );
  INV_X1 U32 ( .A(n65), .ZN(N11) );
  INV_X1 U33 ( .A(n43), .ZN(N31) );
  INV_X1 U34 ( .A(n53), .ZN(N22) );
  INV_X1 U35 ( .A(n52), .ZN(N23) );
  INV_X1 U36 ( .A(n51), .ZN(N24) );
  INV_X1 U37 ( .A(n64), .ZN(N12) );
  INV_X1 U38 ( .A(n63), .ZN(N13) );
  INV_X1 U39 ( .A(n62), .ZN(N14) );
  INV_X1 U40 ( .A(n61), .ZN(N15) );
  INV_X1 U41 ( .A(n60), .ZN(N16) );
  INV_X1 U42 ( .A(n59), .ZN(N17) );
  INV_X1 U43 ( .A(n58), .ZN(N18) );
  INV_X1 U44 ( .A(n57), .ZN(N19) );
  INV_X1 U45 ( .A(n55), .ZN(N20) );
  AOI22_X1 U46 ( .A1(A[2]), .A2(n98), .B1(B[2]), .B2(n101), .ZN(n40) );
  AOI22_X1 U47 ( .A1(A[5]), .A2(n99), .B1(B[5]), .B2(n100), .ZN(n37) );
  AOI22_X1 U48 ( .A1(A[30]), .A2(n99), .B1(B[30]), .B2(n101), .ZN(n42) );
  AOI22_X1 U49 ( .A1(A[6]), .A2(n98), .B1(B[6]), .B2(n100), .ZN(n36) );
  AOI22_X1 U50 ( .A1(A[7]), .A2(n99), .B1(n107), .B2(B[7]), .ZN(n34) );
  AOI22_X1 U51 ( .A1(A[4]), .A2(n98), .B1(B[4]), .B2(n100), .ZN(n38) );
  AOI22_X1 U52 ( .A1(A[31]), .A2(n99), .B1(B[31]), .B2(n101), .ZN(n41) );
  AOI22_X1 U53 ( .A1(A[3]), .A2(n98), .B1(B[3]), .B2(n100), .ZN(n39) );
  AOI22_X1 U54 ( .A1(A[23]), .A2(n98), .B1(B[23]), .B2(n103), .ZN(n50) );
  AOI22_X1 U55 ( .A1(A[1]), .A2(n98), .B1(B[1]), .B2(n102), .ZN(n45) );
  AOI22_X1 U56 ( .A1(A[24]), .A2(n99), .B1(B[24]), .B2(n103), .ZN(n49) );
  AOI22_X1 U57 ( .A1(A[25]), .A2(n99), .B1(B[25]), .B2(n102), .ZN(n48) );
  AOI22_X1 U58 ( .A1(A[27]), .A2(n99), .B1(B[27]), .B2(n102), .ZN(n46) );
  AOI22_X1 U59 ( .A1(A[28]), .A2(n98), .B1(B[28]), .B2(n101), .ZN(n44) );
  AOI22_X1 U60 ( .A1(A[0]), .A2(n98), .B1(B[0]), .B2(n105), .ZN(n56) );
  AOI22_X1 U61 ( .A1(A[10]), .A2(n99), .B1(B[10]), .B2(n107), .ZN(n64) );
  AOI22_X1 U62 ( .A1(A[11]), .A2(n98), .B1(B[11]), .B2(n106), .ZN(n63) );
  AOI22_X1 U63 ( .A1(A[12]), .A2(n99), .B1(B[12]), .B2(n106), .ZN(n62) );
  AOI22_X1 U64 ( .A1(A[13]), .A2(n98), .B1(B[13]), .B2(n106), .ZN(n61) );
  AOI22_X1 U65 ( .A1(A[14]), .A2(n98), .B1(B[14]), .B2(n106), .ZN(n60) );
  AOI22_X1 U66 ( .A1(A[15]), .A2(n99), .B1(B[15]), .B2(n105), .ZN(n59) );
  AOI22_X1 U67 ( .A1(A[16]), .A2(n98), .B1(B[16]), .B2(n105), .ZN(n58) );
  AOI22_X1 U68 ( .A1(A[17]), .A2(n99), .B1(B[17]), .B2(n105), .ZN(n57) );
  AOI22_X1 U69 ( .A1(A[18]), .A2(n99), .B1(B[18]), .B2(n104), .ZN(n55) );
  AOI22_X1 U70 ( .A1(A[19]), .A2(n98), .B1(B[19]), .B2(n104), .ZN(n54) );
  AOI22_X1 U71 ( .A1(A[26]), .A2(n99), .B1(B[26]), .B2(n102), .ZN(n47) );
  AOI22_X1 U72 ( .A1(A[8]), .A2(n98), .B1(B[8]), .B2(n107), .ZN(n66) );
  AOI22_X1 U73 ( .A1(A[9]), .A2(n99), .B1(B[9]), .B2(n107), .ZN(n65) );
  AOI22_X1 U74 ( .A1(A[29]), .A2(n99), .B1(B[29]), .B2(n104), .ZN(n43) );
  AOI22_X1 U75 ( .A1(A[20]), .A2(n99), .B1(B[20]), .B2(n104), .ZN(n53) );
  AOI22_X1 U76 ( .A1(A[21]), .A2(n98), .B1(B[21]), .B2(n103), .ZN(n52) );
  AOI22_X1 U77 ( .A1(A[22]), .A2(n98), .B1(B[22]), .B2(n103), .ZN(n51) );
  INV_X1 U78 ( .A(n108), .ZN(n99) );
endmodule


module compare_N32 ( num1, num2, less, equal, greater );
  input [31:0] num1;
  input [31:0] num2;
  output less, equal, greater;
  wire   n55, n56, n57, n58, n60, n61, n62, n64, n65, n67, n68, n69, n71, n72,
         n74, n75, n76, n77, n80, n81, n82, n83, n86, n87, n88, n89, n90, n92,
         n93, n94, n95, n96, n97, n98, n100, n101, n103, n104, n105, n108,
         n109, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n127, n130, n131, n133, n134, n135,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n151, n152, n153, n154, n155, n157, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335,
         n336, n337, n338, n339, n340, n341;

  NOR3_X2 U4 ( .A1(greater), .A2(n57), .A3(n58), .ZN(equal) );
  NAND3_X1 U106 ( .A1(n81), .A2(n82), .A3(n83), .ZN(n80) );
  NAND3_X1 U107 ( .A1(n87), .A2(n88), .A3(n89), .ZN(n86) );
  NAND3_X1 U108 ( .A1(n135), .A2(n318), .A3(num1[0]), .ZN(n134) );
  NAND3_X1 U109 ( .A1(n82), .A2(n137), .A3(n144), .ZN(n142) );
  NAND3_X1 U110 ( .A1(n94), .A2(n96), .A3(n75), .ZN(n154) );
  NAND2_X1 U2 ( .A1(num2[22]), .A2(n332), .ZN(n83) );
  NOR2_X1 U3 ( .A1(n118), .A2(num1[6]), .ZN(n122) );
  AND2_X1 U5 ( .A1(num1[9]), .A2(n111), .ZN(n300) );
  AND2_X1 U6 ( .A1(num1[8]), .A2(n112), .ZN(n301) );
  NOR3_X1 U7 ( .A1(n300), .A2(n301), .A3(n113), .ZN(n108) );
  NAND2_X1 U8 ( .A1(num1[25]), .A2(n74), .ZN(n302) );
  NAND2_X1 U9 ( .A1(n75), .A2(n76), .ZN(n303) );
  NAND2_X1 U10 ( .A1(num1[24]), .A2(n77), .ZN(n304) );
  AND3_X1 U11 ( .A1(n302), .A2(n303), .A3(n304), .ZN(n71) );
  AND2_X1 U12 ( .A1(n105), .A2(n104), .ZN(n308) );
  NOR2_X1 U13 ( .A1(n308), .A2(n310), .ZN(n100) );
  INV_X1 U14 ( .A(num1[13]), .ZN(n306) );
  NOR2_X1 U15 ( .A1(num2[13]), .A2(n306), .ZN(n307) );
  INV_X1 U16 ( .A(num1[12]), .ZN(n309) );
  NOR2_X1 U17 ( .A1(num2[12]), .A2(n309), .ZN(n305) );
  OR2_X1 U18 ( .A1(n307), .A2(n305), .ZN(n310) );
  AND2_X1 U19 ( .A1(n311), .A2(n312), .ZN(n121) );
  NAND2_X1 U20 ( .A1(n125), .A2(n124), .ZN(n311) );
  NOR2_X1 U21 ( .A1(n315), .A2(n313), .ZN(n312) );
  INV_X1 U22 ( .A(num1[5]), .ZN(n314) );
  NOR2_X1 U23 ( .A1(num2[5]), .A2(n314), .ZN(n315) );
  NOR2_X1 U24 ( .A1(num2[4]), .A2(n153), .ZN(n313) );
  INV_X1 U25 ( .A(n57), .ZN(n55) );
  INV_X1 U26 ( .A(n56), .ZN(n58) );
  NOR4_X1 U27 ( .A1(n145), .A2(n146), .A3(n114), .A4(n147), .ZN(n140) );
  INV_X1 U28 ( .A(n89), .ZN(n146) );
  INV_X1 U29 ( .A(n87), .ZN(n147) );
  OAI221_X1 U30 ( .B1(n320), .B2(n319), .C1(n339), .C2(n61), .A(n124), .ZN(
        n148) );
  NAND4_X1 U31 ( .A1(n138), .A2(n139), .A3(n140), .A4(n141), .ZN(n57) );
  NOR4_X1 U32 ( .A1(n142), .A2(n120), .A3(n143), .A4(n122), .ZN(n141) );
  NOR3_X1 U33 ( .A1(n154), .A2(n72), .A3(n155), .ZN(n138) );
  NOR4_X1 U34 ( .A1(n148), .A2(n101), .A3(n109), .A4(n149), .ZN(n139) );
  INV_X1 U35 ( .A(n115), .ZN(n144) );
  INV_X1 U36 ( .A(n135), .ZN(n143) );
  INV_X1 U37 ( .A(n67), .ZN(n155) );
  INV_X1 U38 ( .A(n104), .ZN(n149) );
  AOI21_X1 U39 ( .B1(n55), .B2(n56), .A(greater), .ZN(less) );
  INV_X1 U40 ( .A(n131), .ZN(n127) );
  OAI21_X1 U41 ( .B1(n320), .B2(n131), .A(n319), .ZN(n130) );
  OAI222_X1 U42 ( .A1(num2[29]), .A2(n338), .B1(n64), .B2(n65), .C1(num2[30]), 
        .C2(n340), .ZN(n62) );
  INV_X1 U43 ( .A(n137), .ZN(n64) );
  OAI222_X1 U44 ( .A1(num2[18]), .A2(n90), .B1(num2[19]), .B2(n329), .C1(n92), 
        .C2(n93), .ZN(n88) );
  INV_X1 U45 ( .A(n94), .ZN(n93) );
  INV_X1 U46 ( .A(num2[17]), .ZN(n95) );
  OAI22_X1 U47 ( .A1(n323), .A2(n152), .B1(num1[13]), .B2(n103), .ZN(n101) );
  INV_X1 U48 ( .A(num2[14]), .ZN(n152) );
  OAI221_X1 U49 ( .B1(num2[20]), .B2(n330), .C1(num2[21]), .C2(n331), .A(n86), 
        .ZN(n81) );
  NOR3_X1 U50 ( .A1(n114), .A2(n115), .A3(n116), .ZN(n113) );
  AOI221_X1 U51 ( .B1(num1[7]), .B2(n117), .C1(num1[6]), .C2(n118), .A(n119), 
        .ZN(n116) );
  NOR3_X1 U52 ( .A1(n120), .A2(n121), .A3(n122), .ZN(n119) );
  OAI22_X1 U53 ( .A1(num1[9]), .A2(n111), .B1(num1[10]), .B2(n151), .ZN(n109)
         );
  INV_X1 U54 ( .A(num2[10]), .ZN(n151) );
  AOI22_X1 U55 ( .A1(n337), .A2(num2[28]), .B1(n336), .B2(num2[27]), .ZN(n67)
         );
  AOI22_X1 U56 ( .A1(n153), .A2(num2[4]), .B1(n316), .B2(num2[3]), .ZN(n124)
         );
  INV_X1 U57 ( .A(num1[4]), .ZN(n153) );
  AOI22_X1 U58 ( .A1(n90), .A2(num2[18]), .B1(n328), .B2(num2[17]), .ZN(n94)
         );
  AOI22_X1 U59 ( .A1(n309), .A2(num2[12]), .B1(n317), .B2(num2[11]), .ZN(n104)
         );
  NOR2_X1 U60 ( .A1(n112), .A2(num1[8]), .ZN(n114) );
  NOR2_X1 U61 ( .A1(n123), .A2(num1[5]), .ZN(n120) );
  NOR2_X1 U62 ( .A1(n117), .A2(num1[7]), .ZN(n115) );
  OAI21_X1 U63 ( .B1(num2[1]), .B2(n133), .A(n134), .ZN(n131) );
  AOI22_X1 U64 ( .A1(n326), .A2(num2[16]), .B1(n325), .B2(num2[15]), .ZN(n96)
         );
  AOI22_X1 U65 ( .A1(n67), .A2(n68), .B1(num1[28]), .B2(n69), .ZN(n65) );
  INV_X1 U66 ( .A(num2[28]), .ZN(n69) );
  OAI222_X1 U67 ( .A1(num2[26]), .A2(n335), .B1(n71), .B2(n72), .C1(num2[27]), 
        .C2(n336), .ZN(n68) );
  AOI22_X1 U68 ( .A1(n334), .A2(num2[24]), .B1(n333), .B2(num2[23]), .ZN(n75)
         );
  INV_X1 U69 ( .A(num1[18]), .ZN(n90) );
  NAND2_X1 U70 ( .A1(num2[31]), .A2(n341), .ZN(n56) );
  NAND2_X1 U71 ( .A1(num2[19]), .A2(n329), .ZN(n89) );
  NAND2_X1 U72 ( .A1(num2[20]), .A2(n330), .ZN(n87) );
  NAND2_X1 U73 ( .A1(num2[29]), .A2(n338), .ZN(n137) );
  OAI22_X1 U74 ( .A1(num1[26]), .A2(n157), .B1(num1[25]), .B2(n74), .ZN(n72)
         );
  INV_X1 U75 ( .A(num2[26]), .ZN(n157) );
  INV_X1 U76 ( .A(num2[6]), .ZN(n118) );
  INV_X1 U77 ( .A(num2[8]), .ZN(n112) );
  NAND2_X1 U78 ( .A1(num2[21]), .A2(n331), .ZN(n82) );
  INV_X1 U79 ( .A(num2[9]), .ZN(n111) );
  INV_X1 U80 ( .A(num2[7]), .ZN(n117) );
  INV_X1 U81 ( .A(num2[30]), .ZN(n61) );
  INV_X1 U82 ( .A(num2[13]), .ZN(n103) );
  INV_X1 U83 ( .A(num2[25]), .ZN(n74) );
  INV_X1 U84 ( .A(num2[5]), .ZN(n123) );
  INV_X1 U85 ( .A(num2[16]), .ZN(n98) );
  INV_X1 U86 ( .A(num2[24]), .ZN(n77) );
  INV_X1 U87 ( .A(num1[3]), .ZN(n316) );
  INV_X1 U88 ( .A(num1[11]), .ZN(n317) );
  INV_X1 U89 ( .A(num1[1]), .ZN(n133) );
  NAND2_X1 U90 ( .A1(num2[1]), .A2(n133), .ZN(n135) );
  OAI21_X1 U91 ( .B1(num2[31]), .B2(n341), .A(n60), .ZN(greater) );
  OAI211_X1 U92 ( .C1(n339), .C2(n61), .A(n62), .B(n56), .ZN(n60) );
  OAI221_X1 U93 ( .B1(num2[22]), .B2(n332), .C1(num2[23]), .C2(n333), .A(n80), 
        .ZN(n76) );
  OAI222_X1 U94 ( .A1(num2[10]), .A2(n322), .B1(n108), .B2(n109), .C1(num2[11]), .C2(n317), .ZN(n105) );
  AOI222_X1 U95 ( .A1(n327), .A2(n95), .B1(n96), .B2(n97), .C1(num1[16]), .C2(
        n98), .ZN(n92) );
  OAI222_X1 U96 ( .A1(num2[14]), .A2(n324), .B1(n100), .B2(n101), .C1(num2[15]), .C2(n325), .ZN(n97) );
  OAI221_X1 U97 ( .B1(n127), .B2(n321), .C1(num2[3]), .C2(n316), .A(n130), 
        .ZN(n125) );
  OAI21_X1 U98 ( .B1(num1[0]), .B2(n318), .A(n83), .ZN(n145) );
  INV_X1 U99 ( .A(num2[0]), .ZN(n318) );
  INV_X1 U100 ( .A(num2[2]), .ZN(n319) );
  INV_X1 U101 ( .A(n321), .ZN(n320) );
  INV_X1 U102 ( .A(num1[2]), .ZN(n321) );
  INV_X1 U103 ( .A(num1[10]), .ZN(n322) );
  INV_X1 U104 ( .A(n324), .ZN(n323) );
  INV_X1 U105 ( .A(num1[14]), .ZN(n324) );
  INV_X1 U111 ( .A(num1[15]), .ZN(n325) );
  INV_X1 U112 ( .A(num1[16]), .ZN(n326) );
  INV_X1 U113 ( .A(n328), .ZN(n327) );
  INV_X1 U114 ( .A(num1[17]), .ZN(n328) );
  INV_X1 U115 ( .A(num1[19]), .ZN(n329) );
  INV_X1 U116 ( .A(num1[20]), .ZN(n330) );
  INV_X1 U117 ( .A(num1[21]), .ZN(n331) );
  INV_X1 U118 ( .A(num1[22]), .ZN(n332) );
  INV_X1 U119 ( .A(num1[23]), .ZN(n333) );
  INV_X1 U120 ( .A(num1[24]), .ZN(n334) );
  INV_X1 U121 ( .A(num1[26]), .ZN(n335) );
  INV_X1 U122 ( .A(num1[27]), .ZN(n336) );
  INV_X1 U123 ( .A(num1[28]), .ZN(n337) );
  INV_X1 U124 ( .A(num1[29]), .ZN(n338) );
  INV_X1 U125 ( .A(n340), .ZN(n339) );
  INV_X1 U126 ( .A(num1[30]), .ZN(n340) );
  INV_X1 U127 ( .A(num1[31]), .ZN(n341) );
endmodule


module p4_adder_N32_N_carry4 ( A, B, Cin, SUM );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input Cin;
  wire   n5, n6;
  wire   [31:0] notb;
  wire   [7:0] carry;
  assign n5 = Cin;

  XOR2_X1 U1 ( .A(n6), .B(B[9]), .Z(notb[9]) );
  XOR2_X1 U2 ( .A(n6), .B(B[8]), .Z(notb[8]) );
  XOR2_X1 U3 ( .A(n6), .B(B[7]), .Z(notb[7]) );
  XOR2_X1 U4 ( .A(n6), .B(B[6]), .Z(notb[6]) );
  XOR2_X1 U5 ( .A(n6), .B(B[5]), .Z(notb[5]) );
  XOR2_X1 U6 ( .A(n6), .B(B[4]), .Z(notb[4]) );
  XOR2_X1 U7 ( .A(n6), .B(B[3]), .Z(notb[3]) );
  XOR2_X1 U8 ( .A(n6), .B(B[31]), .Z(notb[31]) );
  XOR2_X1 U9 ( .A(n6), .B(B[30]), .Z(notb[30]) );
  XOR2_X1 U10 ( .A(n6), .B(B[2]), .Z(notb[2]) );
  XOR2_X1 U11 ( .A(n6), .B(B[29]), .Z(notb[29]) );
  XOR2_X1 U12 ( .A(n6), .B(B[28]), .Z(notb[28]) );
  XOR2_X1 U13 ( .A(n6), .B(B[27]), .Z(notb[27]) );
  XOR2_X1 U14 ( .A(n6), .B(B[26]), .Z(notb[26]) );
  XOR2_X1 U15 ( .A(n6), .B(B[25]), .Z(notb[25]) );
  XOR2_X1 U16 ( .A(n6), .B(B[24]), .Z(notb[24]) );
  XOR2_X1 U17 ( .A(n6), .B(B[23]), .Z(notb[23]) );
  XOR2_X1 U18 ( .A(n6), .B(B[22]), .Z(notb[22]) );
  XOR2_X1 U19 ( .A(n6), .B(B[21]), .Z(notb[21]) );
  XOR2_X1 U20 ( .A(n6), .B(B[20]), .Z(notb[20]) );
  XOR2_X1 U21 ( .A(n6), .B(B[1]), .Z(notb[1]) );
  XOR2_X1 U22 ( .A(n6), .B(B[19]), .Z(notb[19]) );
  XOR2_X1 U23 ( .A(n6), .B(B[18]), .Z(notb[18]) );
  XOR2_X1 U24 ( .A(n6), .B(B[17]), .Z(notb[17]) );
  XOR2_X1 U25 ( .A(n6), .B(B[16]), .Z(notb[16]) );
  XOR2_X1 U26 ( .A(n6), .B(B[15]), .Z(notb[15]) );
  XOR2_X1 U27 ( .A(n6), .B(B[14]), .Z(notb[14]) );
  XOR2_X1 U28 ( .A(n6), .B(B[13]), .Z(notb[13]) );
  XOR2_X1 U29 ( .A(n6), .B(B[12]), .Z(notb[12]) );
  XOR2_X1 U30 ( .A(n6), .B(B[11]), .Z(notb[11]) );
  XOR2_X1 U31 ( .A(n6), .B(B[10]), .Z(notb[10]) );
  XOR2_X1 U32 ( .A(n6), .B(B[0]), .Z(notb[0]) );
  sparse_tree_carry_gen_N5 sparsetree ( .A(A), .B(notb), .C0(n6), .Cout(carry)
         );
  sum_generator_N32_N_carry4 sumgen ( .A(A), .B(notb), .Ci({carry, n6}), .Sum(
        SUM) );
  BUF_X2 U33 ( .A(n5), .Z(n6) );
endmodule


module operatore_logic_REG_SIZE32 ( A, B, OUT_LOGIC_AND, OUT_LOGIC_OR, 
        OUT_LOGIC_XOR );
  input [31:0] A;
  input [31:0] B;
  output [31:0] OUT_LOGIC_AND;
  output [31:0] OUT_LOGIC_OR;
  output [31:0] OUT_LOGIC_XOR;
  wire   n65, n67, n69, n71, n73, n76, n79, n81, n85, n87, n89, n91, n93, n95,
         n97, n99, n101, n103, n106, n107, n109, n110, n111, n113, n115, n117,
         n119, n121, n123, n125, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286;

  XOR2_X1 U129 ( .A(B[9]), .B(A[9]), .Z(OUT_LOGIC_XOR[9]) );
  XOR2_X1 U130 ( .A(B[8]), .B(A[8]), .Z(OUT_LOGIC_XOR[8]) );
  XOR2_X1 U131 ( .A(B[7]), .B(A[7]), .Z(OUT_LOGIC_XOR[7]) );
  XOR2_X1 U132 ( .A(B[6]), .B(A[6]), .Z(OUT_LOGIC_XOR[6]) );
  XOR2_X1 U133 ( .A(B[5]), .B(A[5]), .Z(OUT_LOGIC_XOR[5]) );
  XOR2_X1 U134 ( .A(B[4]), .B(A[4]), .Z(OUT_LOGIC_XOR[4]) );
  XOR2_X1 U135 ( .A(B[3]), .B(A[3]), .Z(OUT_LOGIC_XOR[3]) );
  XOR2_X1 U136 ( .A(B[31]), .B(A[31]), .Z(OUT_LOGIC_XOR[31]) );
  XOR2_X1 U137 ( .A(B[30]), .B(A[30]), .Z(OUT_LOGIC_XOR[30]) );
  XOR2_X1 U138 ( .A(B[2]), .B(A[2]), .Z(OUT_LOGIC_XOR[2]) );
  XOR2_X1 U139 ( .A(B[29]), .B(A[29]), .Z(OUT_LOGIC_XOR[29]) );
  XOR2_X1 U140 ( .A(B[28]), .B(A[28]), .Z(OUT_LOGIC_XOR[28]) );
  XOR2_X1 U141 ( .A(B[27]), .B(A[27]), .Z(OUT_LOGIC_XOR[27]) );
  XOR2_X1 U142 ( .A(B[26]), .B(A[26]), .Z(OUT_LOGIC_XOR[26]) );
  XOR2_X1 U143 ( .A(B[25]), .B(A[25]), .Z(OUT_LOGIC_XOR[25]) );
  XOR2_X1 U144 ( .A(B[24]), .B(A[24]), .Z(OUT_LOGIC_XOR[24]) );
  XOR2_X1 U145 ( .A(B[23]), .B(A[23]), .Z(OUT_LOGIC_XOR[23]) );
  XOR2_X1 U146 ( .A(B[22]), .B(A[22]), .Z(OUT_LOGIC_XOR[22]) );
  XOR2_X1 U147 ( .A(B[21]), .B(A[21]), .Z(OUT_LOGIC_XOR[21]) );
  XOR2_X1 U148 ( .A(B[20]), .B(A[20]), .Z(OUT_LOGIC_XOR[20]) );
  XOR2_X1 U149 ( .A(B[1]), .B(A[1]), .Z(OUT_LOGIC_XOR[1]) );
  XOR2_X1 U150 ( .A(B[19]), .B(A[19]), .Z(OUT_LOGIC_XOR[19]) );
  XOR2_X1 U151 ( .A(B[18]), .B(A[18]), .Z(OUT_LOGIC_XOR[18]) );
  XOR2_X1 U152 ( .A(B[17]), .B(A[17]), .Z(OUT_LOGIC_XOR[17]) );
  XOR2_X1 U153 ( .A(B[16]), .B(A[16]), .Z(OUT_LOGIC_XOR[16]) );
  XOR2_X1 U154 ( .A(B[15]), .B(A[15]), .Z(OUT_LOGIC_XOR[15]) );
  XOR2_X1 U155 ( .A(B[14]), .B(A[14]), .Z(OUT_LOGIC_XOR[14]) );
  XOR2_X1 U156 ( .A(B[13]), .B(A[13]), .Z(OUT_LOGIC_XOR[13]) );
  XOR2_X1 U157 ( .A(B[12]), .B(A[12]), .Z(OUT_LOGIC_XOR[12]) );
  XOR2_X1 U158 ( .A(B[11]), .B(A[11]), .Z(OUT_LOGIC_XOR[11]) );
  XOR2_X1 U159 ( .A(B[10]), .B(A[10]), .Z(OUT_LOGIC_XOR[10]) );
  XOR2_X1 U160 ( .A(B[0]), .B(A[0]), .Z(OUT_LOGIC_XOR[0]) );
  INV_X1 U1 ( .A(A[1]), .ZN(n106) );
  NAND2_X1 U2 ( .A1(n260), .A2(n264), .ZN(OUT_LOGIC_OR[0]) );
  NAND2_X1 U3 ( .A1(n253), .A2(n106), .ZN(OUT_LOGIC_OR[1]) );
  NAND2_X1 U4 ( .A1(n261), .A2(n265), .ZN(OUT_LOGIC_OR[2]) );
  NAND2_X1 U5 ( .A1(n95), .A2(n279), .ZN(OUT_LOGIC_OR[24]) );
  NAND2_X1 U6 ( .A1(n99), .A2(n277), .ZN(OUT_LOGIC_OR[22]) );
  NAND2_X1 U7 ( .A1(n93), .A2(n280), .ZN(OUT_LOGIC_OR[25]) );
  NAND2_X1 U8 ( .A1(n103), .A2(n275), .ZN(OUT_LOGIC_OR[20]) );
  NAND2_X1 U9 ( .A1(n107), .A2(n274), .ZN(OUT_LOGIC_OR[19]) );
  NAND2_X1 U10 ( .A1(n85), .A2(n284), .ZN(OUT_LOGIC_OR[29]) );
  NAND2_X1 U11 ( .A1(n113), .A2(n272), .ZN(OUT_LOGIC_OR[16]) );
  NAND2_X1 U12 ( .A1(n119), .A2(n269), .ZN(OUT_LOGIC_OR[13]) );
  NAND2_X1 U13 ( .A1(n91), .A2(n281), .ZN(OUT_LOGIC_OR[26]) );
  NAND2_X1 U14 ( .A1(n87), .A2(n283), .ZN(OUT_LOGIC_OR[28]) );
  NAND2_X1 U15 ( .A1(n73), .A2(n255), .ZN(OUT_LOGIC_OR[5]) );
  NAND2_X1 U16 ( .A1(n115), .A2(n271), .ZN(OUT_LOGIC_OR[15]) );
  NAND2_X1 U17 ( .A1(n117), .A2(n270), .ZN(OUT_LOGIC_OR[14]) );
  NAND2_X1 U18 ( .A1(n67), .A2(n257), .ZN(OUT_LOGIC_OR[8]) );
  NAND2_X1 U19 ( .A1(n79), .A2(n286), .ZN(OUT_LOGIC_OR[31]) );
  NAND2_X1 U20 ( .A1(n121), .A2(n259), .ZN(OUT_LOGIC_OR[12]) );
  NAND2_X1 U21 ( .A1(n263), .A2(n76), .ZN(OUT_LOGIC_OR[4]) );
  NAND2_X1 U22 ( .A1(n101), .A2(n276), .ZN(OUT_LOGIC_OR[21]) );
  NAND2_X1 U23 ( .A1(n97), .A2(n278), .ZN(OUT_LOGIC_OR[23]) );
  NAND2_X1 U24 ( .A1(n71), .A2(n256), .ZN(OUT_LOGIC_OR[6]) );
  NAND2_X1 U25 ( .A1(n123), .A2(n258), .ZN(OUT_LOGIC_OR[11]) );
  NAND2_X1 U26 ( .A1(n111), .A2(n273), .ZN(OUT_LOGIC_OR[17]) );
  NAND2_X1 U27 ( .A1(n69), .A2(n266), .ZN(OUT_LOGIC_OR[7]) );
  NAND2_X1 U28 ( .A1(n89), .A2(n282), .ZN(OUT_LOGIC_OR[27]) );
  NAND2_X1 U29 ( .A1(n81), .A2(n285), .ZN(OUT_LOGIC_OR[30]) );
  NAND2_X1 U30 ( .A1(n65), .A2(n267), .ZN(OUT_LOGIC_OR[9]) );
  NAND2_X1 U31 ( .A1(n125), .A2(n268), .ZN(OUT_LOGIC_OR[10]) );
  NAND2_X1 U32 ( .A1(n109), .A2(n110), .ZN(OUT_LOGIC_OR[18]) );
  NAND2_X1 U33 ( .A1(n262), .A2(n254), .ZN(OUT_LOGIC_OR[3]) );
  NOR2_X1 U34 ( .A1(n261), .A2(n265), .ZN(OUT_LOGIC_AND[2]) );
  NOR2_X1 U35 ( .A1(n73), .A2(n255), .ZN(OUT_LOGIC_AND[5]) );
  NOR2_X1 U36 ( .A1(n81), .A2(n285), .ZN(OUT_LOGIC_AND[30]) );
  NOR2_X1 U37 ( .A1(n71), .A2(n256), .ZN(OUT_LOGIC_AND[6]) );
  NOR2_X1 U38 ( .A1(n69), .A2(n266), .ZN(OUT_LOGIC_AND[7]) );
  NOR2_X1 U39 ( .A1(n263), .A2(n76), .ZN(OUT_LOGIC_AND[4]) );
  NOR2_X1 U40 ( .A1(n79), .A2(n286), .ZN(OUT_LOGIC_AND[31]) );
  NOR2_X1 U41 ( .A1(n262), .A2(n254), .ZN(OUT_LOGIC_AND[3]) );
  NOR2_X1 U42 ( .A1(n97), .A2(n278), .ZN(OUT_LOGIC_AND[23]) );
  NOR2_X1 U43 ( .A1(n253), .A2(n106), .ZN(OUT_LOGIC_AND[1]) );
  NOR2_X1 U44 ( .A1(n95), .A2(n279), .ZN(OUT_LOGIC_AND[24]) );
  NOR2_X1 U45 ( .A1(n93), .A2(n280), .ZN(OUT_LOGIC_AND[25]) );
  NOR2_X1 U46 ( .A1(n89), .A2(n282), .ZN(OUT_LOGIC_AND[27]) );
  NOR2_X1 U47 ( .A1(n87), .A2(n283), .ZN(OUT_LOGIC_AND[28]) );
  NOR2_X1 U48 ( .A1(n260), .A2(n264), .ZN(OUT_LOGIC_AND[0]) );
  NOR2_X1 U49 ( .A1(n107), .A2(n274), .ZN(OUT_LOGIC_AND[19]) );
  NOR2_X1 U50 ( .A1(n91), .A2(n281), .ZN(OUT_LOGIC_AND[26]) );
  NOR2_X1 U51 ( .A1(n67), .A2(n257), .ZN(OUT_LOGIC_AND[8]) );
  NOR2_X1 U52 ( .A1(n65), .A2(n267), .ZN(OUT_LOGIC_AND[9]) );
  NOR2_X1 U53 ( .A1(n85), .A2(n284), .ZN(OUT_LOGIC_AND[29]) );
  NOR2_X1 U54 ( .A1(n103), .A2(n275), .ZN(OUT_LOGIC_AND[20]) );
  NOR2_X1 U55 ( .A1(n101), .A2(n276), .ZN(OUT_LOGIC_AND[21]) );
  NOR2_X1 U56 ( .A1(n99), .A2(n277), .ZN(OUT_LOGIC_AND[22]) );
  NOR2_X1 U57 ( .A1(n125), .A2(n268), .ZN(OUT_LOGIC_AND[10]) );
  NOR2_X1 U58 ( .A1(n123), .A2(n258), .ZN(OUT_LOGIC_AND[11]) );
  NOR2_X1 U59 ( .A1(n121), .A2(n259), .ZN(OUT_LOGIC_AND[12]) );
  NOR2_X1 U60 ( .A1(n119), .A2(n269), .ZN(OUT_LOGIC_AND[13]) );
  NOR2_X1 U61 ( .A1(n117), .A2(n270), .ZN(OUT_LOGIC_AND[14]) );
  NOR2_X1 U62 ( .A1(n115), .A2(n271), .ZN(OUT_LOGIC_AND[15]) );
  NOR2_X1 U63 ( .A1(n113), .A2(n272), .ZN(OUT_LOGIC_AND[16]) );
  NOR2_X1 U64 ( .A1(n111), .A2(n273), .ZN(OUT_LOGIC_AND[17]) );
  NOR2_X1 U65 ( .A1(n109), .A2(n110), .ZN(OUT_LOGIC_AND[18]) );
  INV_X1 U66 ( .A(A[4]), .ZN(n76) );
  INV_X1 U67 ( .A(A[18]), .ZN(n110) );
  INV_X1 U68 ( .A(B[27]), .ZN(n89) );
  INV_X1 U69 ( .A(B[12]), .ZN(n121) );
  INV_X1 U70 ( .A(B[16]), .ZN(n113) );
  INV_X1 U71 ( .A(B[24]), .ZN(n95) );
  INV_X1 U72 ( .A(B[28]), .ZN(n87) );
  INV_X1 U73 ( .A(B[18]), .ZN(n109) );
  INV_X1 U74 ( .A(B[17]), .ZN(n111) );
  INV_X1 U75 ( .A(B[30]), .ZN(n81) );
  INV_X1 U76 ( .A(B[20]), .ZN(n103) );
  INV_X1 U77 ( .A(B[26]), .ZN(n91) );
  INV_X1 U78 ( .A(B[19]), .ZN(n107) );
  INV_X1 U79 ( .A(B[29]), .ZN(n85) );
  INV_X1 U80 ( .A(B[21]), .ZN(n101) );
  INV_X1 U81 ( .A(B[31]), .ZN(n79) );
  INV_X1 U82 ( .A(B[11]), .ZN(n123) );
  INV_X1 U83 ( .A(B[15]), .ZN(n115) );
  INV_X1 U84 ( .A(B[23]), .ZN(n97) );
  INV_X1 U85 ( .A(B[10]), .ZN(n125) );
  INV_X1 U86 ( .A(B[14]), .ZN(n117) );
  INV_X1 U87 ( .A(B[22]), .ZN(n99) );
  INV_X1 U88 ( .A(B[5]), .ZN(n73) );
  INV_X1 U89 ( .A(B[6]), .ZN(n71) );
  INV_X1 U90 ( .A(B[7]), .ZN(n69) );
  INV_X1 U91 ( .A(B[8]), .ZN(n67) );
  INV_X1 U92 ( .A(B[9]), .ZN(n65) );
  INV_X1 U93 ( .A(B[13]), .ZN(n119) );
  INV_X1 U94 ( .A(B[25]), .ZN(n93) );
  INV_X1 U95 ( .A(B[1]), .ZN(n253) );
  INV_X1 U96 ( .A(A[3]), .ZN(n254) );
  INV_X1 U97 ( .A(A[5]), .ZN(n255) );
  INV_X1 U98 ( .A(A[6]), .ZN(n256) );
  INV_X1 U99 ( .A(A[8]), .ZN(n257) );
  INV_X1 U100 ( .A(A[11]), .ZN(n258) );
  INV_X1 U101 ( .A(A[12]), .ZN(n259) );
  INV_X1 U102 ( .A(B[0]), .ZN(n260) );
  INV_X1 U103 ( .A(B[2]), .ZN(n261) );
  INV_X1 U104 ( .A(B[3]), .ZN(n262) );
  INV_X1 U105 ( .A(B[4]), .ZN(n263) );
  INV_X1 U106 ( .A(A[0]), .ZN(n264) );
  INV_X1 U107 ( .A(A[2]), .ZN(n265) );
  INV_X1 U108 ( .A(A[7]), .ZN(n266) );
  INV_X1 U109 ( .A(A[9]), .ZN(n267) );
  INV_X1 U110 ( .A(A[10]), .ZN(n268) );
  INV_X1 U111 ( .A(A[13]), .ZN(n269) );
  INV_X1 U112 ( .A(A[14]), .ZN(n270) );
  INV_X1 U113 ( .A(A[15]), .ZN(n271) );
  INV_X1 U114 ( .A(A[16]), .ZN(n272) );
  INV_X1 U115 ( .A(A[17]), .ZN(n273) );
  INV_X1 U116 ( .A(A[19]), .ZN(n274) );
  INV_X1 U117 ( .A(A[20]), .ZN(n275) );
  INV_X1 U118 ( .A(A[21]), .ZN(n276) );
  INV_X1 U119 ( .A(A[22]), .ZN(n277) );
  INV_X1 U120 ( .A(A[23]), .ZN(n278) );
  INV_X1 U121 ( .A(A[24]), .ZN(n279) );
  INV_X1 U122 ( .A(A[25]), .ZN(n280) );
  INV_X1 U123 ( .A(A[26]), .ZN(n281) );
  INV_X1 U124 ( .A(A[27]), .ZN(n282) );
  INV_X1 U125 ( .A(A[28]), .ZN(n283) );
  INV_X1 U126 ( .A(A[29]), .ZN(n284) );
  INV_X1 U127 ( .A(A[30]), .ZN(n285) );
  INV_X1 U128 ( .A(A[31]), .ZN(n286) );
endmodule


module SHIFTER_GENERIC_N32 ( A, B, LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE, 
        OUTPUT );
  input [31:0] A;
  input [4:0] B;
  output [31:0] OUTPUT;
  input LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE;
  wire   N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N105, N106, N107, N108, N109,
         N110, N111, N112, N113, N114, N115, N116, N117, N118, N119, N120,
         N121, N122, N123, N124, N125, N126, N127, N128, N129, N130, N131,
         N132, N133, N134, N135, N136, N137, N138, N139, N140, N141, N142,
         N143, N144, N145, N146, N147, N148, N149, N150, N151, N152, N153,
         N154, N155, N156, N157, N158, N159, N160, N161, N162, N163, N164,
         N165, N166, N167, N168, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N224, N225, N226, N227, N228, N229, N230,
         N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, N241,
         N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252,
         N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263,
         N264, N265, n171, n192, n193, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213;
  assign n171 = B[1];
  assign n192 = B[3];
  assign n193 = B[4];

  SHIFTER_GENERIC_N32_DW01_ash_0 C88 ( .A(A), .DATA_TC(1'b0), .SH({n213, n212, 
        B[2], n171, B[0]}), .SH_TC(1'b0), .B({N265, N264, N263, N262, N261, 
        N260, N259, N258, N257, N256, N255, N254, N253, N252, N251, N250, N249, 
        N248, N247, N246, N245, N244, N243, N242, N241, N240, N239, N238, N237, 
        N236, N235, N234}) );
  SHIFTER_GENERIC_N32_DW_sla_0 C86 ( .A(A), .SH({n213, n212, B[2], n171, B[0]}), .SH_TC(1'b0), .B({N233, N232, N231, N230, N229, N228, N227, N226, N225, N224, 
        N223, N222, N221, N220, N219, N218, N217, N216, N215, N214, N213, N212, 
        N211, N210, N209, N208, N207, N206, N205, N204, N203, N202}) );
  SHIFTER_GENERIC_N32_DW_rash_0 C50 ( .A(A), .DATA_TC(1'b0), .SH({n213, n212, 
        B[2], n171, B[0]}), .SH_TC(1'b0), .B({N168, N167, N166, N165, N164, 
        N163, N162, N161, N160, N159, N158, N157, N156, N155, N154, N153, N152, 
        N151, N150, N149, N148, N147, N146, N145, N144, N143, N142, N141, N140, 
        N139, N138, N137}) );
  SHIFTER_GENERIC_N32_DW_sra_0 C48 ( .A(A), .SH({n213, n212, B[2], n171, B[0]}), .SH_TC(1'b0), .B({N136, N135, N134, N133, N132, N131, N130, N129, N128, N127, 
        N126, N125, N124, N123, N122, N121, N120, N119, N118, N117, N116, N115, 
        N114, N113, N112, N111, N110, N109, N108, N107, N106, N105}) );
  SHIFTER_GENERIC_N32_DW_lbsh_0 C10 ( .A(A), .SH({n213, n212, B[2], n171, B[0]}), .SH_TC(1'b0), .B({N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, 
        N59, N58, N57, N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, 
        N45, N44, N43, N42, N41, N40, N39}) );
  SHIFTER_GENERIC_N32_DW_rbsh_0 C8 ( .A(A), .SH({n213, n212, B[2], n171, B[0]}), .SH_TC(1'b0), .B({N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7}) );
  BUF_X1 U5 ( .A(n192), .Z(n212) );
  NAND2_X1 U6 ( .A1(n27), .A2(n28), .ZN(OUTPUT[6]) );
  AOI222_X1 U7 ( .A1(N45), .A2(n202), .B1(N13), .B2(n199), .C1(N240), .C2(n196), .ZN(n27) );
  AOI222_X1 U8 ( .A1(N208), .A2(n211), .B1(N143), .B2(n208), .C1(N111), .C2(
        n205), .ZN(n28) );
  NAND2_X1 U9 ( .A1(n25), .A2(n26), .ZN(OUTPUT[7]) );
  AOI222_X1 U10 ( .A1(N46), .A2(n202), .B1(N14), .B2(n199), .C1(N241), .C2(
        n196), .ZN(n25) );
  AOI222_X1 U13 ( .A1(N209), .A2(n211), .B1(N144), .B2(n208), .C1(N112), .C2(
        n205), .ZN(n26) );
  NAND2_X1 U14 ( .A1(n23), .A2(n24), .ZN(OUTPUT[8]) );
  AOI222_X1 U15 ( .A1(N47), .A2(n202), .B1(N15), .B2(n199), .C1(N242), .C2(
        n196), .ZN(n23) );
  AOI222_X1 U16 ( .A1(N210), .A2(n211), .B1(N145), .B2(n208), .C1(N113), .C2(
        n205), .ZN(n24) );
  NAND2_X1 U17 ( .A1(n15), .A2(n16), .ZN(OUTPUT[9]) );
  AOI222_X1 U18 ( .A1(N48), .A2(n202), .B1(N16), .B2(n199), .C1(N243), .C2(
        n196), .ZN(n15) );
  AOI222_X1 U19 ( .A1(N211), .A2(n211), .B1(N146), .B2(n208), .C1(N114), .C2(
        n205), .ZN(n16) );
  NAND2_X1 U20 ( .A1(n83), .A2(n84), .ZN(OUTPUT[0]) );
  AOI222_X1 U21 ( .A1(N39), .A2(n200), .B1(N7), .B2(n197), .C1(N234), .C2(n194), .ZN(n83) );
  AOI222_X1 U22 ( .A1(N202), .A2(n209), .B1(N137), .B2(n206), .C1(N105), .C2(
        n203), .ZN(n84) );
  NAND2_X1 U23 ( .A1(n61), .A2(n62), .ZN(OUTPUT[1]) );
  AOI222_X1 U24 ( .A1(N40), .A2(n201), .B1(N8), .B2(n197), .C1(N235), .C2(n194), .ZN(n61) );
  AOI222_X1 U25 ( .A1(N203), .A2(n210), .B1(N138), .B2(n206), .C1(N106), .C2(
        n203), .ZN(n62) );
  NAND2_X1 U26 ( .A1(n81), .A2(n82), .ZN(OUTPUT[10]) );
  AOI222_X1 U27 ( .A1(N49), .A2(n200), .B1(N17), .B2(n197), .C1(N244), .C2(
        n194), .ZN(n81) );
  AOI222_X1 U28 ( .A1(N212), .A2(n209), .B1(N147), .B2(n206), .C1(N115), .C2(
        n203), .ZN(n82) );
  NAND2_X1 U29 ( .A1(n79), .A2(n80), .ZN(OUTPUT[11]) );
  AOI222_X1 U30 ( .A1(N50), .A2(n200), .B1(N18), .B2(n197), .C1(N245), .C2(
        n194), .ZN(n79) );
  AOI222_X1 U31 ( .A1(N213), .A2(n209), .B1(N148), .B2(n206), .C1(N116), .C2(
        n203), .ZN(n80) );
  NAND2_X1 U32 ( .A1(n77), .A2(n78), .ZN(OUTPUT[12]) );
  AOI222_X1 U33 ( .A1(N51), .A2(n200), .B1(N19), .B2(n197), .C1(N246), .C2(
        n194), .ZN(n77) );
  AOI222_X1 U34 ( .A1(N214), .A2(n209), .B1(N149), .B2(n206), .C1(N117), .C2(
        n203), .ZN(n78) );
  NAND2_X1 U35 ( .A1(n75), .A2(n76), .ZN(OUTPUT[13]) );
  AOI222_X1 U36 ( .A1(N52), .A2(n200), .B1(N20), .B2(n197), .C1(N247), .C2(
        n194), .ZN(n75) );
  AOI222_X1 U37 ( .A1(N215), .A2(n209), .B1(N150), .B2(n206), .C1(N118), .C2(
        n203), .ZN(n76) );
  NAND2_X1 U38 ( .A1(n73), .A2(n74), .ZN(OUTPUT[14]) );
  AOI222_X1 U39 ( .A1(N53), .A2(n200), .B1(N21), .B2(n197), .C1(N248), .C2(
        n194), .ZN(n73) );
  AOI222_X1 U40 ( .A1(N216), .A2(n209), .B1(N151), .B2(n206), .C1(N119), .C2(
        n203), .ZN(n74) );
  NAND2_X1 U41 ( .A1(n71), .A2(n72), .ZN(OUTPUT[15]) );
  AOI222_X1 U42 ( .A1(N54), .A2(n200), .B1(N22), .B2(n197), .C1(N249), .C2(
        n194), .ZN(n71) );
  AOI222_X1 U43 ( .A1(N217), .A2(n209), .B1(N152), .B2(n206), .C1(N120), .C2(
        n203), .ZN(n72) );
  NAND2_X1 U44 ( .A1(n69), .A2(n70), .ZN(OUTPUT[16]) );
  AOI222_X1 U45 ( .A1(N55), .A2(n200), .B1(N23), .B2(n197), .C1(N250), .C2(
        n194), .ZN(n69) );
  AOI222_X1 U46 ( .A1(N218), .A2(n209), .B1(N153), .B2(n206), .C1(N121), .C2(
        n203), .ZN(n70) );
  NAND2_X1 U47 ( .A1(n67), .A2(n68), .ZN(OUTPUT[17]) );
  AOI222_X1 U48 ( .A1(N56), .A2(n200), .B1(N24), .B2(n197), .C1(N251), .C2(
        n194), .ZN(n67) );
  AOI222_X1 U49 ( .A1(N219), .A2(n209), .B1(N154), .B2(n206), .C1(N122), .C2(
        n203), .ZN(n68) );
  NAND2_X1 U50 ( .A1(n65), .A2(n66), .ZN(OUTPUT[18]) );
  AOI222_X1 U51 ( .A1(N57), .A2(n200), .B1(N25), .B2(n197), .C1(N252), .C2(
        n194), .ZN(n65) );
  AOI222_X1 U52 ( .A1(N220), .A2(n209), .B1(N155), .B2(n206), .C1(N123), .C2(
        n203), .ZN(n66) );
  NAND2_X1 U53 ( .A1(n63), .A2(n64), .ZN(OUTPUT[19]) );
  AOI222_X1 U54 ( .A1(N58), .A2(n200), .B1(N26), .B2(n197), .C1(N253), .C2(
        n194), .ZN(n63) );
  AOI222_X1 U55 ( .A1(N221), .A2(n209), .B1(N156), .B2(n206), .C1(N124), .C2(
        n203), .ZN(n64) );
  NAND2_X1 U56 ( .A1(n59), .A2(n60), .ZN(OUTPUT[20]) );
  AOI222_X1 U57 ( .A1(N59), .A2(n201), .B1(N27), .B2(n198), .C1(N254), .C2(
        n195), .ZN(n59) );
  AOI222_X1 U58 ( .A1(N222), .A2(n210), .B1(N157), .B2(n207), .C1(N125), .C2(
        n204), .ZN(n60) );
  NAND2_X1 U59 ( .A1(n57), .A2(n58), .ZN(OUTPUT[21]) );
  AOI222_X1 U60 ( .A1(N60), .A2(n201), .B1(N28), .B2(n198), .C1(N255), .C2(
        n195), .ZN(n57) );
  AOI222_X1 U61 ( .A1(N223), .A2(n210), .B1(N158), .B2(n207), .C1(N126), .C2(
        n204), .ZN(n58) );
  NAND2_X1 U62 ( .A1(n55), .A2(n56), .ZN(OUTPUT[22]) );
  AOI222_X1 U63 ( .A1(N61), .A2(n201), .B1(N29), .B2(n198), .C1(N256), .C2(
        n195), .ZN(n55) );
  AOI222_X1 U64 ( .A1(N224), .A2(n210), .B1(N159), .B2(n207), .C1(N127), .C2(
        n204), .ZN(n56) );
  NAND2_X1 U65 ( .A1(n53), .A2(n54), .ZN(OUTPUT[23]) );
  AOI222_X1 U66 ( .A1(N62), .A2(n201), .B1(N30), .B2(n198), .C1(N257), .C2(
        n195), .ZN(n53) );
  AOI222_X1 U67 ( .A1(N225), .A2(n210), .B1(N160), .B2(n207), .C1(N128), .C2(
        n204), .ZN(n54) );
  NAND2_X1 U68 ( .A1(n51), .A2(n52), .ZN(OUTPUT[24]) );
  AOI222_X1 U69 ( .A1(N63), .A2(n201), .B1(N31), .B2(n198), .C1(N258), .C2(
        n195), .ZN(n51) );
  AOI222_X1 U70 ( .A1(N226), .A2(n210), .B1(N161), .B2(n207), .C1(N129), .C2(
        n204), .ZN(n52) );
  NAND2_X1 U71 ( .A1(n49), .A2(n50), .ZN(OUTPUT[25]) );
  AOI222_X1 U72 ( .A1(N64), .A2(n201), .B1(N32), .B2(n198), .C1(N259), .C2(
        n195), .ZN(n49) );
  AOI222_X1 U73 ( .A1(N227), .A2(n210), .B1(N162), .B2(n207), .C1(N130), .C2(
        n204), .ZN(n50) );
  NAND2_X1 U74 ( .A1(n47), .A2(n48), .ZN(OUTPUT[26]) );
  AOI222_X1 U75 ( .A1(N65), .A2(n201), .B1(N33), .B2(n198), .C1(N260), .C2(
        n195), .ZN(n47) );
  AOI222_X1 U76 ( .A1(N228), .A2(n210), .B1(N163), .B2(n207), .C1(N131), .C2(
        n204), .ZN(n48) );
  NAND2_X1 U77 ( .A1(n45), .A2(n46), .ZN(OUTPUT[27]) );
  AOI222_X1 U78 ( .A1(N66), .A2(n201), .B1(N34), .B2(n198), .C1(N261), .C2(
        n195), .ZN(n45) );
  AOI222_X1 U79 ( .A1(N229), .A2(n210), .B1(N164), .B2(n207), .C1(N132), .C2(
        n204), .ZN(n46) );
  NAND2_X1 U80 ( .A1(n31), .A2(n32), .ZN(OUTPUT[4]) );
  AOI222_X1 U81 ( .A1(N43), .A2(n202), .B1(N11), .B2(n199), .C1(N238), .C2(
        n196), .ZN(n31) );
  AOI222_X1 U82 ( .A1(N206), .A2(n211), .B1(N141), .B2(n208), .C1(N109), .C2(
        n205), .ZN(n32) );
  NAND2_X1 U83 ( .A1(n29), .A2(n30), .ZN(OUTPUT[5]) );
  AOI222_X1 U84 ( .A1(N44), .A2(n202), .B1(N12), .B2(n199), .C1(N239), .C2(
        n196), .ZN(n29) );
  AOI222_X1 U85 ( .A1(N207), .A2(n211), .B1(N142), .B2(n208), .C1(N110), .C2(
        n205), .ZN(n30) );
  BUF_X1 U86 ( .A(n20), .Z(n200) );
  BUF_X1 U87 ( .A(n20), .Z(n201) );
  BUF_X1 U88 ( .A(n20), .Z(n202) );
  BUF_X1 U89 ( .A(n18), .Z(n206) );
  BUF_X1 U90 ( .A(n18), .Z(n207) );
  BUF_X1 U91 ( .A(n19), .Z(n203) );
  BUF_X1 U92 ( .A(n19), .Z(n204) );
  BUF_X1 U93 ( .A(n18), .Z(n208) );
  BUF_X1 U94 ( .A(n19), .Z(n205) );
  NAND2_X1 U95 ( .A1(n33), .A2(n34), .ZN(OUTPUT[3]) );
  AOI222_X1 U96 ( .A1(N42), .A2(n202), .B1(N10), .B2(n199), .C1(N237), .C2(
        n196), .ZN(n33) );
  AOI222_X1 U97 ( .A1(N205), .A2(n211), .B1(N140), .B2(n208), .C1(N108), .C2(
        n205), .ZN(n34) );
  NAND2_X1 U98 ( .A1(n39), .A2(n40), .ZN(OUTPUT[2]) );
  AOI222_X1 U99 ( .A1(N41), .A2(n202), .B1(N9), .B2(n198), .C1(N236), .C2(n195), .ZN(n39) );
  AOI222_X1 U100 ( .A1(N204), .A2(n211), .B1(N139), .B2(n207), .C1(N107), .C2(
        n204), .ZN(n40) );
  NAND2_X1 U101 ( .A1(n43), .A2(n44), .ZN(OUTPUT[28]) );
  AOI222_X1 U102 ( .A1(N67), .A2(n201), .B1(N35), .B2(n198), .C1(N262), .C2(
        n195), .ZN(n43) );
  AOI222_X1 U103 ( .A1(N230), .A2(n210), .B1(N165), .B2(n207), .C1(N133), .C2(
        n204), .ZN(n44) );
  NAND2_X1 U104 ( .A1(n41), .A2(n42), .ZN(OUTPUT[29]) );
  AOI222_X1 U105 ( .A1(N68), .A2(n201), .B1(N36), .B2(n198), .C1(N263), .C2(
        n195), .ZN(n41) );
  AOI222_X1 U106 ( .A1(N231), .A2(n210), .B1(N166), .B2(n207), .C1(N134), .C2(
        n204), .ZN(n42) );
  NAND2_X1 U107 ( .A1(n37), .A2(n38), .ZN(OUTPUT[30]) );
  AOI222_X1 U108 ( .A1(N69), .A2(n202), .B1(N37), .B2(n198), .C1(N264), .C2(
        n195), .ZN(n37) );
  AOI222_X1 U109 ( .A1(N232), .A2(n211), .B1(N167), .B2(n207), .C1(N135), .C2(
        n204), .ZN(n38) );
  NAND2_X1 U110 ( .A1(n35), .A2(n36), .ZN(OUTPUT[31]) );
  AOI222_X1 U111 ( .A1(N70), .A2(n202), .B1(N38), .B2(n199), .C1(N265), .C2(
        n196), .ZN(n35) );
  AOI222_X1 U112 ( .A1(N233), .A2(n211), .B1(N168), .B2(n208), .C1(N136), .C2(
        n205), .ZN(n36) );
  BUF_X1 U113 ( .A(n21), .Z(n197) );
  BUF_X1 U114 ( .A(n21), .Z(n198) );
  BUF_X1 U115 ( .A(n17), .Z(n209) );
  BUF_X1 U116 ( .A(n17), .Z(n210) );
  BUF_X1 U117 ( .A(n17), .Z(n211) );
  BUF_X1 U118 ( .A(n22), .Z(n194) );
  BUF_X1 U119 ( .A(n22), .Z(n195) );
  BUF_X1 U120 ( .A(n21), .Z(n199) );
  BUF_X1 U121 ( .A(n22), .Z(n196) );
  NOR2_X1 U122 ( .A1(n85), .A2(SHIFT_ROTATE), .ZN(n20) );
  AND3_X1 U123 ( .A1(LOGIC_ARITH), .A2(n85), .A3(SHIFT_ROTATE), .ZN(n18) );
  AND3_X1 U124 ( .A1(n85), .A2(n86), .A3(SHIFT_ROTATE), .ZN(n19) );
  INV_X1 U125 ( .A(LOGIC_ARITH), .ZN(n86) );
  CLKBUF_X1 U126 ( .A(n193), .Z(n213) );
  NOR2_X1 U127 ( .A1(LEFT_RIGHT), .A2(SHIFT_ROTATE), .ZN(n21) );
  AND3_X1 U128 ( .A1(SHIFT_ROTATE), .A2(LOGIC_ARITH), .A3(LEFT_RIGHT), .ZN(n22) );
  INV_X1 U129 ( .A(LEFT_RIGHT), .ZN(n85) );
  AND3_X1 U130 ( .A1(SHIFT_ROTATE), .A2(n86), .A3(LEFT_RIGHT), .ZN(n17) );
endmodule


module RCA_GEN_NBIT32 ( A, B, Ci, S, Co );
  input [31:0] A;
  input [31:0] B;
  output [31:0] S;
  input Ci;
  output Co;

  wire   [31:1] CTMP;

  FA_0 fai_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_95 fai_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_94 fai_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_93 fai_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(CTMP[4]) );
  FA_92 fai_5 ( .A(A[4]), .B(B[4]), .Ci(CTMP[4]), .S(S[4]), .Co(CTMP[5]) );
  FA_91 fai_6 ( .A(A[5]), .B(B[5]), .Ci(CTMP[5]), .S(S[5]), .Co(CTMP[6]) );
  FA_90 fai_7 ( .A(A[6]), .B(B[6]), .Ci(CTMP[6]), .S(S[6]), .Co(CTMP[7]) );
  FA_89 fai_8 ( .A(A[7]), .B(B[7]), .Ci(CTMP[7]), .S(S[7]), .Co(CTMP[8]) );
  FA_88 fai_9 ( .A(A[8]), .B(B[8]), .Ci(CTMP[8]), .S(S[8]), .Co(CTMP[9]) );
  FA_87 fai_10 ( .A(A[9]), .B(B[9]), .Ci(CTMP[9]), .S(S[9]), .Co(CTMP[10]) );
  FA_86 fai_11 ( .A(A[10]), .B(B[10]), .Ci(CTMP[10]), .S(S[10]), .Co(CTMP[11])
         );
  FA_85 fai_12 ( .A(A[11]), .B(B[11]), .Ci(CTMP[11]), .S(S[11]), .Co(CTMP[12])
         );
  FA_84 fai_13 ( .A(A[12]), .B(B[12]), .Ci(CTMP[12]), .S(S[12]), .Co(CTMP[13])
         );
  FA_83 fai_14 ( .A(A[13]), .B(B[13]), .Ci(CTMP[13]), .S(S[13]), .Co(CTMP[14])
         );
  FA_82 fai_15 ( .A(A[14]), .B(B[14]), .Ci(CTMP[14]), .S(S[14]), .Co(CTMP[15])
         );
  FA_81 fai_16 ( .A(A[15]), .B(B[15]), .Ci(CTMP[15]), .S(S[15]), .Co(CTMP[16])
         );
  FA_80 fai_17 ( .A(A[16]), .B(B[16]), .Ci(CTMP[16]), .S(S[16]), .Co(CTMP[17])
         );
  FA_79 fai_18 ( .A(A[17]), .B(B[17]), .Ci(CTMP[17]), .S(S[17]), .Co(CTMP[18])
         );
  FA_78 fai_19 ( .A(A[18]), .B(B[18]), .Ci(CTMP[18]), .S(S[18]), .Co(CTMP[19])
         );
  FA_77 fai_20 ( .A(A[19]), .B(B[19]), .Ci(CTMP[19]), .S(S[19]), .Co(CTMP[20])
         );
  FA_76 fai_21 ( .A(A[20]), .B(B[20]), .Ci(CTMP[20]), .S(S[20]), .Co(CTMP[21])
         );
  FA_75 fai_22 ( .A(A[21]), .B(B[21]), .Ci(CTMP[21]), .S(S[21]), .Co(CTMP[22])
         );
  FA_74 fai_23 ( .A(A[22]), .B(B[22]), .Ci(CTMP[22]), .S(S[22]), .Co(CTMP[23])
         );
  FA_73 fai_24 ( .A(A[23]), .B(B[23]), .Ci(CTMP[23]), .S(S[23]), .Co(CTMP[24])
         );
  FA_72 fai_25 ( .A(A[24]), .B(B[24]), .Ci(CTMP[24]), .S(S[24]), .Co(CTMP[25])
         );
  FA_71 fai_26 ( .A(A[25]), .B(B[25]), .Ci(CTMP[25]), .S(S[25]), .Co(CTMP[26])
         );
  FA_70 fai_27 ( .A(A[26]), .B(B[26]), .Ci(CTMP[26]), .S(S[26]), .Co(CTMP[27])
         );
  FA_69 fai_28 ( .A(A[27]), .B(B[27]), .Ci(CTMP[27]), .S(S[27]), .Co(CTMP[28])
         );
  FA_68 fai_29 ( .A(A[28]), .B(B[28]), .Ci(CTMP[28]), .S(S[28]), .Co(CTMP[29])
         );
  FA_67 fai_30 ( .A(A[29]), .B(B[29]), .Ci(CTMP[29]), .S(S[29]), .Co(CTMP[30])
         );
  FA_66 fai_31 ( .A(A[30]), .B(B[30]), .Ci(CTMP[30]), .S(S[30]), .Co(CTMP[31])
         );
  FA_65 fai_32 ( .A(A[31]), .B(B[31]), .Ci(CTMP[31]), .S(S[31]), .Co(Co) );
endmodule


module mux21_N5 ( A, B, SEL, Y );
  input [4:0] A;
  input [4:0] B;
  output [4:0] Y;
  input SEL;
  wire   n7, n8, n9, n10, n11, n12;

  INV_X1 U1 ( .A(SEL), .ZN(n8) );
  INV_X1 U2 ( .A(n10), .ZN(Y[2]) );
  AOI22_X1 U3 ( .A1(A[2]), .A2(n8), .B1(B[2]), .B2(SEL), .ZN(n10) );
  INV_X1 U4 ( .A(n11), .ZN(Y[1]) );
  AOI22_X1 U5 ( .A1(A[1]), .A2(n8), .B1(B[1]), .B2(SEL), .ZN(n11) );
  INV_X1 U6 ( .A(n12), .ZN(Y[0]) );
  AOI22_X1 U7 ( .A1(A[0]), .A2(n8), .B1(B[0]), .B2(SEL), .ZN(n12) );
  INV_X1 U8 ( .A(n7), .ZN(Y[4]) );
  AOI22_X1 U9 ( .A1(A[4]), .A2(n8), .B1(SEL), .B2(B[4]), .ZN(n7) );
  INV_X1 U10 ( .A(n9), .ZN(Y[3]) );
  AOI22_X1 U11 ( .A1(A[3]), .A2(n8), .B1(B[3]), .B2(SEL), .ZN(n9) );
endmodule


module mux21_N32_1 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136;

  INV_X1 U1 ( .A(n136), .ZN(n126) );
  INV_X1 U2 ( .A(n136), .ZN(n127) );
  BUF_X1 U3 ( .A(n123), .Z(n128) );
  BUF_X1 U4 ( .A(n125), .Z(n134) );
  BUF_X1 U5 ( .A(n124), .Z(n133) );
  BUF_X1 U6 ( .A(n124), .Z(n131) );
  BUF_X1 U7 ( .A(n123), .Z(n130) );
  BUF_X1 U8 ( .A(n124), .Z(n132) );
  BUF_X1 U9 ( .A(n123), .Z(n129) );
  BUF_X1 U10 ( .A(n125), .Z(n136) );
  BUF_X1 U11 ( .A(n125), .Z(n135) );
  INV_X1 U12 ( .A(n42), .ZN(Y[31]) );
  AOI22_X1 U13 ( .A1(A[31]), .A2(n126), .B1(B[31]), .B2(n129), .ZN(n42) );
  INV_X1 U14 ( .A(n66), .ZN(Y[0]) );
  AOI22_X1 U15 ( .A1(A[0]), .A2(n126), .B1(B[0]), .B2(n135), .ZN(n66) );
  INV_X1 U16 ( .A(n55), .ZN(Y[1]) );
  AOI22_X1 U17 ( .A1(A[1]), .A2(n126), .B1(B[1]), .B2(n132), .ZN(n55) );
  INV_X1 U18 ( .A(n44), .ZN(Y[2]) );
  AOI22_X1 U19 ( .A1(A[2]), .A2(n127), .B1(B[2]), .B2(n129), .ZN(n44) );
  INV_X1 U20 ( .A(n41), .ZN(Y[3]) );
  AOI22_X1 U21 ( .A1(A[3]), .A2(n127), .B1(B[3]), .B2(n129), .ZN(n41) );
  INV_X1 U22 ( .A(n40), .ZN(Y[4]) );
  AOI22_X1 U23 ( .A1(A[4]), .A2(n126), .B1(B[4]), .B2(n129), .ZN(n40) );
  INV_X1 U24 ( .A(n39), .ZN(Y[5]) );
  AOI22_X1 U25 ( .A1(A[5]), .A2(n127), .B1(B[5]), .B2(n128), .ZN(n39) );
  INV_X1 U26 ( .A(n38), .ZN(Y[6]) );
  AOI22_X1 U27 ( .A1(A[6]), .A2(n126), .B1(B[6]), .B2(n128), .ZN(n38) );
  INV_X1 U28 ( .A(n37), .ZN(Y[7]) );
  AOI22_X1 U29 ( .A1(A[7]), .A2(n127), .B1(B[7]), .B2(n128), .ZN(n37) );
  INV_X1 U30 ( .A(n36), .ZN(Y[8]) );
  AOI22_X1 U31 ( .A1(A[8]), .A2(n126), .B1(B[8]), .B2(n128), .ZN(n36) );
  INV_X1 U32 ( .A(n34), .ZN(Y[9]) );
  AOI22_X1 U33 ( .A1(A[9]), .A2(n127), .B1(n135), .B2(B[9]), .ZN(n34) );
  INV_X1 U34 ( .A(n65), .ZN(Y[10]) );
  AOI22_X1 U35 ( .A1(A[10]), .A2(n126), .B1(B[10]), .B2(n135), .ZN(n65) );
  INV_X1 U36 ( .A(n64), .ZN(Y[11]) );
  AOI22_X1 U37 ( .A1(A[11]), .A2(n126), .B1(B[11]), .B2(n135), .ZN(n64) );
  INV_X1 U38 ( .A(n63), .ZN(Y[12]) );
  AOI22_X1 U39 ( .A1(A[12]), .A2(n126), .B1(B[12]), .B2(n134), .ZN(n63) );
  INV_X1 U40 ( .A(n62), .ZN(Y[13]) );
  AOI22_X1 U41 ( .A1(A[13]), .A2(n126), .B1(B[13]), .B2(n134), .ZN(n62) );
  INV_X1 U42 ( .A(n61), .ZN(Y[14]) );
  AOI22_X1 U43 ( .A1(A[14]), .A2(n126), .B1(B[14]), .B2(n134), .ZN(n61) );
  INV_X1 U44 ( .A(n60), .ZN(Y[15]) );
  AOI22_X1 U45 ( .A1(A[15]), .A2(n126), .B1(B[15]), .B2(n134), .ZN(n60) );
  INV_X1 U46 ( .A(n59), .ZN(Y[16]) );
  AOI22_X1 U47 ( .A1(A[16]), .A2(n126), .B1(B[16]), .B2(n133), .ZN(n59) );
  INV_X1 U48 ( .A(n58), .ZN(Y[17]) );
  AOI22_X1 U49 ( .A1(A[17]), .A2(n126), .B1(B[17]), .B2(n133), .ZN(n58) );
  INV_X1 U50 ( .A(n57), .ZN(Y[18]) );
  AOI22_X1 U51 ( .A1(A[18]), .A2(n126), .B1(B[18]), .B2(n133), .ZN(n57) );
  INV_X1 U52 ( .A(n56), .ZN(Y[19]) );
  AOI22_X1 U53 ( .A1(A[19]), .A2(n126), .B1(B[19]), .B2(n133), .ZN(n56) );
  INV_X1 U54 ( .A(n54), .ZN(Y[20]) );
  AOI22_X1 U55 ( .A1(A[20]), .A2(n127), .B1(B[20]), .B2(n132), .ZN(n54) );
  INV_X1 U56 ( .A(n53), .ZN(Y[21]) );
  AOI22_X1 U57 ( .A1(A[21]), .A2(n127), .B1(B[21]), .B2(n132), .ZN(n53) );
  INV_X1 U58 ( .A(n52), .ZN(Y[22]) );
  AOI22_X1 U59 ( .A1(A[22]), .A2(n127), .B1(B[22]), .B2(n131), .ZN(n52) );
  INV_X1 U60 ( .A(n51), .ZN(Y[23]) );
  AOI22_X1 U61 ( .A1(A[23]), .A2(n127), .B1(B[23]), .B2(n131), .ZN(n51) );
  INV_X1 U62 ( .A(n50), .ZN(Y[24]) );
  AOI22_X1 U63 ( .A1(A[24]), .A2(n127), .B1(B[24]), .B2(n131), .ZN(n50) );
  INV_X1 U64 ( .A(n49), .ZN(Y[25]) );
  AOI22_X1 U65 ( .A1(A[25]), .A2(n127), .B1(B[25]), .B2(n131), .ZN(n49) );
  INV_X1 U66 ( .A(n48), .ZN(Y[26]) );
  AOI22_X1 U67 ( .A1(A[26]), .A2(n127), .B1(B[26]), .B2(n130), .ZN(n48) );
  INV_X1 U68 ( .A(n47), .ZN(Y[27]) );
  AOI22_X1 U69 ( .A1(A[27]), .A2(n127), .B1(B[27]), .B2(n130), .ZN(n47) );
  INV_X1 U70 ( .A(n46), .ZN(Y[28]) );
  AOI22_X1 U71 ( .A1(A[28]), .A2(n127), .B1(B[28]), .B2(n130), .ZN(n46) );
  INV_X1 U72 ( .A(n45), .ZN(Y[29]) );
  AOI22_X1 U73 ( .A1(A[29]), .A2(n127), .B1(B[29]), .B2(n130), .ZN(n45) );
  INV_X1 U74 ( .A(n43), .ZN(Y[30]) );
  AOI22_X1 U75 ( .A1(A[30]), .A2(n127), .B1(B[30]), .B2(n132), .ZN(n43) );
  BUF_X1 U76 ( .A(SEL), .Z(n125) );
  BUF_X1 U77 ( .A(SEL), .Z(n124) );
  BUF_X1 U78 ( .A(SEL), .Z(n123) );
endmodule


module registro_N5_1 ( data, enable, clock, clear, Q );
  input [4:0] data;
  output [4:0] Q;
  input enable, clock, clear;
  wire   n1, n2, n3, n4, n5, net44880, net44881, net44882, net44883, net44884,
         n6, n7, n8, n9, n10;

  DFFR_X1 \Q_reg[4]  ( .D(n1), .CK(clock), .RN(clear), .Q(Q[4]), .QN(net44884)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n2), .CK(clock), .RN(clear), .Q(Q[3]), .QN(net44883)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n3), .CK(clock), .RN(clear), .Q(Q[2]), .QN(net44882)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n4), .CK(clock), .RN(clear), .Q(Q[1]), .QN(net44881)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n5), .CK(clock), .RN(clear), .Q(Q[0]), .QN(net44880)
         );
  OAI21_X1 U2 ( .B1(net44880), .B2(enable), .A(n6), .ZN(n5) );
  NAND2_X1 U3 ( .A1(enable), .A2(data[0]), .ZN(n6) );
  OAI21_X1 U4 ( .B1(net44881), .B2(enable), .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(enable), .ZN(n7) );
  OAI21_X1 U6 ( .B1(net44882), .B2(enable), .A(n8), .ZN(n3) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(enable), .ZN(n8) );
  OAI21_X1 U8 ( .B1(net44883), .B2(enable), .A(n9), .ZN(n2) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(enable), .ZN(n9) );
  OAI21_X1 U10 ( .B1(net44884), .B2(enable), .A(n10), .ZN(n1) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(enable), .ZN(n10) );
endmodule


module registro_N32_1 ( data, enable, clock, clear, Q );
  input [31:0] data;
  output [31:0] Q;
  input enable, clock, clear;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net44624, net44625, net44626, net44627, net44628, net44629,
         net44630, net44631, net44632, net44633, net44634, net44635, net44636,
         net44637, net44638, net44639, net44640, net44641, net44642, net44643,
         net44644, net44645, net44646, net44647, net44648, net44649, net44650,
         net44651, net44652, net44653, net44654, net44655, n167, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n174, n175, n176, n177, n178, n179, n180, n181, n182;
  assign n167 = clear;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(clock), .RN(n176), .Q(Q[31]), .QN(net44655) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(clock), .RN(n176), .Q(Q[30]), .QN(net44654) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(clock), .RN(n176), .Q(Q[29]), .QN(net44653) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(clock), .RN(n176), .Q(Q[28]), .QN(net44652) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(clock), .RN(n176), .Q(Q[27]), .QN(net44651) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(clock), .RN(n176), .Q(Q[26]), .QN(net44650) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(clock), .RN(n176), .Q(Q[25]), .QN(net44649) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(clock), .RN(n176), .Q(Q[24]), .QN(net44648) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(clock), .RN(n176), .Q(Q[23]), .QN(net44647) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(clock), .RN(n176), .Q(Q[22]), .QN(
        net44646) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(clock), .RN(n174), .Q(Q[21]), .QN(
        net44645) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(clock), .RN(n174), .Q(Q[20]), .QN(
        net44644) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(clock), .RN(n174), .Q(Q[19]), .QN(
        net44643) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(clock), .RN(n174), .Q(Q[18]), .QN(
        net44642) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(clock), .RN(n174), .Q(Q[17]), .QN(
        net44641) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(clock), .RN(n174), .Q(Q[16]), .QN(
        net44640) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(clock), .RN(n174), .Q(Q[15]), .QN(
        net44639) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(clock), .RN(n174), .Q(Q[14]), .QN(
        net44638) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(clock), .RN(n174), .Q(Q[13]), .QN(
        net44637) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(clock), .RN(n174), .Q(Q[12]), .QN(
        net44636) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(clock), .RN(n174), .Q(Q[11]), .QN(
        net44635) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(clock), .RN(n175), .Q(Q[10]), .QN(
        net44634) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(clock), .RN(n175), .Q(Q[9]), .QN(net44633)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(clock), .RN(n175), .Q(Q[8]), .QN(net44632)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(clock), .RN(n175), .Q(Q[7]), .QN(net44631)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(clock), .RN(n175), .Q(Q[6]), .QN(net44630)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(clock), .RN(n175), .Q(Q[5]), .QN(net44629)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(clock), .RN(n175), .Q(Q[4]), .QN(net44628)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(clock), .RN(n175), .Q(Q[3]), .QN(net44627)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(clock), .RN(n175), .Q(Q[2]), .QN(net44626)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(clock), .RN(n175), .Q(Q[1]), .QN(net44625)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(clock), .RN(n175), .Q(Q[0]), .QN(net44624)
         );
  BUF_X1 U2 ( .A(n167), .Z(n175) );
  BUF_X1 U3 ( .A(n167), .Z(n174) );
  BUF_X1 U4 ( .A(n167), .Z(n176) );
  BUF_X1 U5 ( .A(enable), .Z(n178) );
  BUF_X1 U6 ( .A(enable), .Z(n177) );
  BUF_X1 U7 ( .A(enable), .Z(n179) );
  BUF_X1 U8 ( .A(enable), .Z(n181) );
  BUF_X1 U9 ( .A(enable), .Z(n180) );
  OAI21_X1 U10 ( .B1(net44625), .B2(n179), .A(n40), .ZN(n31) );
  NAND2_X1 U11 ( .A1(data[1]), .A2(n178), .ZN(n40) );
  OAI21_X1 U12 ( .B1(net44648), .B2(n179), .A(n34), .ZN(n8) );
  NAND2_X1 U13 ( .A1(data[24]), .A2(n177), .ZN(n34) );
  OAI21_X1 U14 ( .B1(net44649), .B2(n179), .A(n35), .ZN(n7) );
  NAND2_X1 U15 ( .A1(data[25]), .A2(n177), .ZN(n35) );
  OAI21_X1 U16 ( .B1(net44651), .B2(n179), .A(n37), .ZN(n5) );
  NAND2_X1 U17 ( .A1(data[27]), .A2(n177), .ZN(n37) );
  OAI21_X1 U18 ( .B1(net44652), .B2(n179), .A(n38), .ZN(n4) );
  NAND2_X1 U19 ( .A1(data[28]), .A2(n178), .ZN(n38) );
  OAI21_X1 U20 ( .B1(net44624), .B2(n180), .A(n39), .ZN(n32) );
  NAND2_X1 U21 ( .A1(data[0]), .A2(n178), .ZN(n39) );
  OAI21_X1 U22 ( .B1(net44626), .B2(n180), .A(n41), .ZN(n30) );
  NAND2_X1 U23 ( .A1(data[2]), .A2(n178), .ZN(n41) );
  OAI21_X1 U24 ( .B1(net44627), .B2(n180), .A(n43), .ZN(n29) );
  NAND2_X1 U25 ( .A1(data[3]), .A2(n178), .ZN(n43) );
  OAI21_X1 U26 ( .B1(net44628), .B2(n180), .A(n44), .ZN(n28) );
  NAND2_X1 U27 ( .A1(data[4]), .A2(n179), .ZN(n44) );
  OAI21_X1 U28 ( .B1(net44629), .B2(n180), .A(n45), .ZN(n27) );
  NAND2_X1 U29 ( .A1(data[5]), .A2(n179), .ZN(n45) );
  OAI21_X1 U30 ( .B1(net44630), .B2(n180), .A(n46), .ZN(n26) );
  NAND2_X1 U31 ( .A1(data[6]), .A2(n179), .ZN(n46) );
  OAI21_X1 U32 ( .B1(net44631), .B2(n180), .A(n47), .ZN(n25) );
  NAND2_X1 U33 ( .A1(data[7]), .A2(n179), .ZN(n47) );
  OAI21_X1 U34 ( .B1(net44632), .B2(n180), .A(n48), .ZN(n24) );
  NAND2_X1 U35 ( .A1(data[8]), .A2(n179), .ZN(n48) );
  OAI21_X1 U36 ( .B1(net44633), .B2(n181), .A(n49), .ZN(n23) );
  NAND2_X1 U37 ( .A1(data[9]), .A2(n179), .ZN(n49) );
  OAI21_X1 U38 ( .B1(net44634), .B2(n181), .A(n50), .ZN(n22) );
  NAND2_X1 U39 ( .A1(data[10]), .A2(n178), .ZN(n50) );
  OAI21_X1 U40 ( .B1(net44635), .B2(n181), .A(n51), .ZN(n21) );
  NAND2_X1 U41 ( .A1(data[11]), .A2(n178), .ZN(n51) );
  OAI21_X1 U42 ( .B1(net44636), .B2(n181), .A(n52), .ZN(n20) );
  NAND2_X1 U43 ( .A1(data[12]), .A2(n178), .ZN(n52) );
  OAI21_X1 U44 ( .B1(net44637), .B2(n181), .A(n54), .ZN(n19) );
  NAND2_X1 U45 ( .A1(data[13]), .A2(n178), .ZN(n54) );
  OAI21_X1 U46 ( .B1(net44638), .B2(n181), .A(n55), .ZN(n18) );
  NAND2_X1 U47 ( .A1(data[14]), .A2(n178), .ZN(n55) );
  OAI21_X1 U48 ( .B1(net44639), .B2(n181), .A(n56), .ZN(n17) );
  NAND2_X1 U49 ( .A1(data[15]), .A2(n178), .ZN(n56) );
  OAI21_X1 U50 ( .B1(net44640), .B2(n181), .A(n57), .ZN(n16) );
  NAND2_X1 U51 ( .A1(data[16]), .A2(n177), .ZN(n57) );
  OAI21_X1 U52 ( .B1(net44641), .B2(n181), .A(n58), .ZN(n15) );
  NAND2_X1 U53 ( .A1(data[17]), .A2(n177), .ZN(n58) );
  OAI21_X1 U54 ( .B1(net44642), .B2(n181), .A(n59), .ZN(n14) );
  NAND2_X1 U55 ( .A1(data[18]), .A2(n177), .ZN(n59) );
  OAI21_X1 U56 ( .B1(net44643), .B2(n181), .A(n60), .ZN(n13) );
  NAND2_X1 U57 ( .A1(data[19]), .A2(n177), .ZN(n60) );
  OAI21_X1 U58 ( .B1(net44647), .B2(n180), .A(n33), .ZN(n9) );
  NAND2_X1 U59 ( .A1(n182), .A2(data[23]), .ZN(n33) );
  OAI21_X1 U60 ( .B1(net44650), .B2(n180), .A(n36), .ZN(n6) );
  NAND2_X1 U61 ( .A1(data[26]), .A2(n177), .ZN(n36) );
  OAI21_X1 U62 ( .B1(net44653), .B2(n180), .A(n42), .ZN(n3) );
  NAND2_X1 U63 ( .A1(data[29]), .A2(n179), .ZN(n42) );
  OAI21_X1 U64 ( .B1(net44654), .B2(n181), .A(n53), .ZN(n2) );
  NAND2_X1 U65 ( .A1(data[30]), .A2(n178), .ZN(n53) );
  OAI21_X1 U66 ( .B1(net44655), .B2(n180), .A(n64), .ZN(n1) );
  NAND2_X1 U67 ( .A1(data[31]), .A2(n177), .ZN(n64) );
  OAI21_X1 U68 ( .B1(net44644), .B2(n182), .A(n61), .ZN(n12) );
  NAND2_X1 U69 ( .A1(data[20]), .A2(n177), .ZN(n61) );
  OAI21_X1 U70 ( .B1(net44645), .B2(n182), .A(n62), .ZN(n11) );
  NAND2_X1 U71 ( .A1(data[21]), .A2(n177), .ZN(n62) );
  OAI21_X1 U72 ( .B1(net44646), .B2(n182), .A(n63), .ZN(n10) );
  NAND2_X1 U73 ( .A1(data[22]), .A2(n177), .ZN(n63) );
  CLKBUF_X1 U74 ( .A(enable), .Z(n182) );
endmodule


module registro_N32_2 ( data, enable, clock, clear, Q );
  input [31:0] data;
  output [31:0] Q;
  input enable, clock, clear;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net44624, net44625, net44626, net44627, net44628, net44629,
         net44630, net44631, net44632, net44633, net44634, net44635, net44636,
         net44637, net44638, net44639, net44640, net44641, net44642, net44643,
         net44644, net44645, net44646, net44647, net44648, net44649, net44650,
         net44651, net44652, net44653, net44654, net44655, n135, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n142, n143, n144, n145, n146, n147, n148, n149, n150;
  assign n135 = clear;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(clock), .RN(n144), .Q(Q[31]), .QN(net44655) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(clock), .RN(n144), .Q(Q[30]), .QN(net44654) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(clock), .RN(n144), .Q(Q[29]), .QN(net44653) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(clock), .RN(n144), .Q(Q[28]), .QN(net44652) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(clock), .RN(n144), .Q(Q[27]), .QN(net44651) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(clock), .RN(n144), .Q(Q[26]), .QN(net44650) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(clock), .RN(n144), .Q(Q[25]), .QN(net44649) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(clock), .RN(n144), .Q(Q[24]), .QN(net44648) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(clock), .RN(n144), .Q(Q[23]), .QN(net44647) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(clock), .RN(n144), .Q(Q[22]), .QN(
        net44646) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(clock), .RN(n142), .Q(Q[21]), .QN(
        net44645) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(clock), .RN(n142), .Q(Q[20]), .QN(
        net44644) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(clock), .RN(n142), .Q(Q[19]), .QN(
        net44643) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(clock), .RN(n142), .Q(Q[18]), .QN(
        net44642) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(clock), .RN(n142), .Q(Q[17]), .QN(
        net44641) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(clock), .RN(n142), .Q(Q[16]), .QN(
        net44640) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(clock), .RN(n142), .Q(Q[15]), .QN(
        net44639) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(clock), .RN(n142), .Q(Q[14]), .QN(
        net44638) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(clock), .RN(n142), .Q(Q[13]), .QN(
        net44637) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(clock), .RN(n142), .Q(Q[12]), .QN(
        net44636) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(clock), .RN(n142), .Q(Q[11]), .QN(
        net44635) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(clock), .RN(n143), .Q(Q[10]), .QN(
        net44634) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(clock), .RN(n143), .Q(Q[9]), .QN(net44633)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(clock), .RN(n143), .Q(Q[8]), .QN(net44632)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(clock), .RN(n143), .Q(Q[7]), .QN(net44631)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(clock), .RN(n143), .Q(Q[6]), .QN(net44630)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(clock), .RN(n143), .Q(Q[5]), .QN(net44629)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(clock), .RN(n143), .Q(Q[4]), .QN(net44628)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(clock), .RN(n143), .Q(Q[3]), .QN(net44627)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(clock), .RN(n143), .Q(Q[2]), .QN(net44626)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(clock), .RN(n143), .Q(Q[1]), .QN(net44625)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(clock), .RN(n143), .Q(Q[0]), .QN(net44624)
         );
  BUF_X1 U2 ( .A(n135), .Z(n143) );
  BUF_X1 U3 ( .A(n135), .Z(n142) );
  BUF_X1 U4 ( .A(n135), .Z(n144) );
  OAI21_X1 U5 ( .B1(net44624), .B2(n148), .A(n39), .ZN(n32) );
  NAND2_X1 U6 ( .A1(data[0]), .A2(n146), .ZN(n39) );
  OAI21_X1 U7 ( .B1(net44625), .B2(n147), .A(n40), .ZN(n31) );
  NAND2_X1 U8 ( .A1(data[1]), .A2(n146), .ZN(n40) );
  OAI21_X1 U9 ( .B1(net44626), .B2(n148), .A(n41), .ZN(n30) );
  NAND2_X1 U10 ( .A1(data[2]), .A2(n146), .ZN(n41) );
  OAI21_X1 U11 ( .B1(net44634), .B2(n149), .A(n50), .ZN(n22) );
  NAND2_X1 U12 ( .A1(data[10]), .A2(n146), .ZN(n50) );
  OAI21_X1 U13 ( .B1(net44635), .B2(n149), .A(n51), .ZN(n21) );
  NAND2_X1 U14 ( .A1(data[11]), .A2(n146), .ZN(n51) );
  OAI21_X1 U15 ( .B1(net44636), .B2(n149), .A(n52), .ZN(n20) );
  NAND2_X1 U16 ( .A1(data[12]), .A2(n146), .ZN(n52) );
  OAI21_X1 U17 ( .B1(net44637), .B2(n149), .A(n54), .ZN(n19) );
  NAND2_X1 U18 ( .A1(data[13]), .A2(n146), .ZN(n54) );
  OAI21_X1 U19 ( .B1(net44638), .B2(n149), .A(n55), .ZN(n18) );
  NAND2_X1 U20 ( .A1(data[14]), .A2(n146), .ZN(n55) );
  OAI21_X1 U21 ( .B1(net44639), .B2(n149), .A(n56), .ZN(n17) );
  NAND2_X1 U22 ( .A1(data[15]), .A2(n146), .ZN(n56) );
  OAI21_X1 U23 ( .B1(net44640), .B2(n149), .A(n57), .ZN(n16) );
  NAND2_X1 U24 ( .A1(data[16]), .A2(n145), .ZN(n57) );
  OAI21_X1 U25 ( .B1(net44641), .B2(n149), .A(n58), .ZN(n15) );
  NAND2_X1 U26 ( .A1(data[17]), .A2(n145), .ZN(n58) );
  OAI21_X1 U27 ( .B1(net44642), .B2(n149), .A(n59), .ZN(n14) );
  NAND2_X1 U28 ( .A1(data[18]), .A2(n145), .ZN(n59) );
  OAI21_X1 U29 ( .B1(net44643), .B2(n149), .A(n60), .ZN(n13) );
  NAND2_X1 U30 ( .A1(data[19]), .A2(n145), .ZN(n60) );
  OAI21_X1 U31 ( .B1(net44644), .B2(n150), .A(n61), .ZN(n12) );
  NAND2_X1 U32 ( .A1(data[20]), .A2(n145), .ZN(n61) );
  OAI21_X1 U33 ( .B1(net44645), .B2(n150), .A(n62), .ZN(n11) );
  NAND2_X1 U34 ( .A1(data[21]), .A2(n145), .ZN(n62) );
  OAI21_X1 U35 ( .B1(net44646), .B2(n150), .A(n63), .ZN(n10) );
  NAND2_X1 U36 ( .A1(data[22]), .A2(n145), .ZN(n63) );
  OAI21_X1 U37 ( .B1(net44648), .B2(n147), .A(n34), .ZN(n8) );
  NAND2_X1 U38 ( .A1(data[24]), .A2(n145), .ZN(n34) );
  OAI21_X1 U39 ( .B1(net44649), .B2(n147), .A(n35), .ZN(n7) );
  NAND2_X1 U40 ( .A1(data[25]), .A2(n145), .ZN(n35) );
  OAI21_X1 U41 ( .B1(net44650), .B2(n148), .A(n36), .ZN(n6) );
  NAND2_X1 U42 ( .A1(data[26]), .A2(n145), .ZN(n36) );
  OAI21_X1 U43 ( .B1(net44651), .B2(n147), .A(n37), .ZN(n5) );
  NAND2_X1 U44 ( .A1(data[27]), .A2(n145), .ZN(n37) );
  OAI21_X1 U45 ( .B1(net44652), .B2(n147), .A(n38), .ZN(n4) );
  NAND2_X1 U46 ( .A1(data[28]), .A2(n146), .ZN(n38) );
  OAI21_X1 U47 ( .B1(net44654), .B2(n149), .A(n53), .ZN(n2) );
  NAND2_X1 U48 ( .A1(data[30]), .A2(n146), .ZN(n53) );
  OAI21_X1 U49 ( .B1(net44653), .B2(n148), .A(n42), .ZN(n3) );
  NAND2_X1 U50 ( .A1(data[29]), .A2(n147), .ZN(n42) );
  OAI21_X1 U51 ( .B1(net44647), .B2(n148), .A(n33), .ZN(n9) );
  NAND2_X1 U52 ( .A1(n150), .A2(data[23]), .ZN(n33) );
  OAI21_X1 U53 ( .B1(net44627), .B2(n148), .A(n43), .ZN(n29) );
  NAND2_X1 U54 ( .A1(data[3]), .A2(n146), .ZN(n43) );
  OAI21_X1 U55 ( .B1(net44628), .B2(n148), .A(n44), .ZN(n28) );
  NAND2_X1 U56 ( .A1(data[4]), .A2(n147), .ZN(n44) );
  OAI21_X1 U57 ( .B1(net44629), .B2(n148), .A(n45), .ZN(n27) );
  NAND2_X1 U58 ( .A1(data[5]), .A2(n147), .ZN(n45) );
  OAI21_X1 U59 ( .B1(net44630), .B2(n148), .A(n46), .ZN(n26) );
  NAND2_X1 U60 ( .A1(data[6]), .A2(n147), .ZN(n46) );
  OAI21_X1 U61 ( .B1(net44631), .B2(n148), .A(n47), .ZN(n25) );
  NAND2_X1 U62 ( .A1(data[7]), .A2(n147), .ZN(n47) );
  OAI21_X1 U63 ( .B1(net44632), .B2(n148), .A(n48), .ZN(n24) );
  NAND2_X1 U64 ( .A1(data[8]), .A2(n147), .ZN(n48) );
  OAI21_X1 U65 ( .B1(net44633), .B2(n149), .A(n49), .ZN(n23) );
  NAND2_X1 U66 ( .A1(data[9]), .A2(n147), .ZN(n49) );
  OAI21_X1 U67 ( .B1(net44655), .B2(n148), .A(n64), .ZN(n1) );
  NAND2_X1 U68 ( .A1(data[31]), .A2(n145), .ZN(n64) );
  BUF_X1 U69 ( .A(enable), .Z(n146) );
  BUF_X1 U70 ( .A(enable), .Z(n145) );
  BUF_X1 U71 ( .A(enable), .Z(n147) );
  BUF_X1 U72 ( .A(enable), .Z(n149) );
  BUF_X1 U73 ( .A(enable), .Z(n148) );
  CLKBUF_X1 U74 ( .A(enable), .Z(n150) );
endmodule


module mux21_N32_2 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n123, n124, n125, n126, n127, n128, n129, n130,
         n131, n132, n133, n134, n135, n136;

  INV_X1 U1 ( .A(n136), .ZN(n126) );
  INV_X1 U2 ( .A(n136), .ZN(n127) );
  BUF_X1 U3 ( .A(n125), .Z(n136) );
  BUF_X1 U4 ( .A(n123), .Z(n128) );
  BUF_X1 U5 ( .A(n125), .Z(n134) );
  BUF_X1 U6 ( .A(n124), .Z(n133) );
  BUF_X1 U7 ( .A(n124), .Z(n131) );
  BUF_X1 U8 ( .A(n123), .Z(n130) );
  BUF_X1 U9 ( .A(n124), .Z(n132) );
  BUF_X1 U10 ( .A(n123), .Z(n129) );
  BUF_X1 U11 ( .A(n125), .Z(n135) );
  INV_X1 U12 ( .A(n66), .ZN(Y[0]) );
  AOI22_X1 U13 ( .A1(A[0]), .A2(n126), .B1(B[0]), .B2(n135), .ZN(n66) );
  INV_X1 U14 ( .A(n55), .ZN(Y[1]) );
  AOI22_X1 U15 ( .A1(A[1]), .A2(n126), .B1(B[1]), .B2(n132), .ZN(n55) );
  INV_X1 U16 ( .A(n44), .ZN(Y[2]) );
  AOI22_X1 U17 ( .A1(A[2]), .A2(n127), .B1(B[2]), .B2(n129), .ZN(n44) );
  INV_X1 U18 ( .A(n65), .ZN(Y[10]) );
  AOI22_X1 U19 ( .A1(A[10]), .A2(n126), .B1(B[10]), .B2(n135), .ZN(n65) );
  INV_X1 U20 ( .A(n64), .ZN(Y[11]) );
  AOI22_X1 U21 ( .A1(A[11]), .A2(n126), .B1(B[11]), .B2(n135), .ZN(n64) );
  INV_X1 U22 ( .A(n63), .ZN(Y[12]) );
  AOI22_X1 U23 ( .A1(A[12]), .A2(n126), .B1(B[12]), .B2(n134), .ZN(n63) );
  INV_X1 U24 ( .A(n62), .ZN(Y[13]) );
  AOI22_X1 U25 ( .A1(A[13]), .A2(n126), .B1(B[13]), .B2(n134), .ZN(n62) );
  INV_X1 U26 ( .A(n61), .ZN(Y[14]) );
  AOI22_X1 U27 ( .A1(A[14]), .A2(n126), .B1(B[14]), .B2(n134), .ZN(n61) );
  INV_X1 U28 ( .A(n60), .ZN(Y[15]) );
  AOI22_X1 U29 ( .A1(A[15]), .A2(n126), .B1(B[15]), .B2(n134), .ZN(n60) );
  INV_X1 U30 ( .A(n59), .ZN(Y[16]) );
  AOI22_X1 U31 ( .A1(A[16]), .A2(n126), .B1(B[16]), .B2(n133), .ZN(n59) );
  INV_X1 U32 ( .A(n58), .ZN(Y[17]) );
  AOI22_X1 U33 ( .A1(A[17]), .A2(n126), .B1(B[17]), .B2(n133), .ZN(n58) );
  INV_X1 U34 ( .A(n57), .ZN(Y[18]) );
  AOI22_X1 U35 ( .A1(A[18]), .A2(n126), .B1(B[18]), .B2(n133), .ZN(n57) );
  INV_X1 U36 ( .A(n56), .ZN(Y[19]) );
  AOI22_X1 U37 ( .A1(A[19]), .A2(n126), .B1(B[19]), .B2(n133), .ZN(n56) );
  INV_X1 U38 ( .A(n54), .ZN(Y[20]) );
  AOI22_X1 U39 ( .A1(A[20]), .A2(n127), .B1(B[20]), .B2(n132), .ZN(n54) );
  INV_X1 U40 ( .A(n53), .ZN(Y[21]) );
  AOI22_X1 U41 ( .A1(A[21]), .A2(n127), .B1(B[21]), .B2(n132), .ZN(n53) );
  INV_X1 U42 ( .A(n52), .ZN(Y[22]) );
  AOI22_X1 U43 ( .A1(A[22]), .A2(n127), .B1(B[22]), .B2(n131), .ZN(n52) );
  INV_X1 U44 ( .A(n50), .ZN(Y[24]) );
  AOI22_X1 U45 ( .A1(A[24]), .A2(n127), .B1(B[24]), .B2(n131), .ZN(n50) );
  INV_X1 U46 ( .A(n49), .ZN(Y[25]) );
  AOI22_X1 U47 ( .A1(A[25]), .A2(n127), .B1(B[25]), .B2(n131), .ZN(n49) );
  INV_X1 U48 ( .A(n48), .ZN(Y[26]) );
  AOI22_X1 U49 ( .A1(A[26]), .A2(n127), .B1(B[26]), .B2(n130), .ZN(n48) );
  INV_X1 U50 ( .A(n47), .ZN(Y[27]) );
  AOI22_X1 U51 ( .A1(A[27]), .A2(n127), .B1(B[27]), .B2(n130), .ZN(n47) );
  INV_X1 U52 ( .A(n46), .ZN(Y[28]) );
  AOI22_X1 U53 ( .A1(A[28]), .A2(n127), .B1(B[28]), .B2(n130), .ZN(n46) );
  INV_X1 U54 ( .A(n43), .ZN(Y[30]) );
  AOI22_X1 U55 ( .A1(A[30]), .A2(n127), .B1(B[30]), .B2(n132), .ZN(n43) );
  INV_X1 U56 ( .A(n45), .ZN(Y[29]) );
  AOI22_X1 U57 ( .A1(A[29]), .A2(n127), .B1(B[29]), .B2(n130), .ZN(n45) );
  INV_X1 U58 ( .A(n51), .ZN(Y[23]) );
  AOI22_X1 U59 ( .A1(A[23]), .A2(n127), .B1(B[23]), .B2(n131), .ZN(n51) );
  INV_X1 U60 ( .A(n41), .ZN(Y[3]) );
  AOI22_X1 U61 ( .A1(A[3]), .A2(n126), .B1(B[3]), .B2(n129), .ZN(n41) );
  INV_X1 U62 ( .A(n40), .ZN(Y[4]) );
  AOI22_X1 U63 ( .A1(A[4]), .A2(n127), .B1(B[4]), .B2(n129), .ZN(n40) );
  INV_X1 U64 ( .A(n39), .ZN(Y[5]) );
  AOI22_X1 U65 ( .A1(A[5]), .A2(n126), .B1(B[5]), .B2(n128), .ZN(n39) );
  INV_X1 U66 ( .A(n38), .ZN(Y[6]) );
  AOI22_X1 U67 ( .A1(A[6]), .A2(n127), .B1(B[6]), .B2(n128), .ZN(n38) );
  INV_X1 U68 ( .A(n37), .ZN(Y[7]) );
  AOI22_X1 U69 ( .A1(A[7]), .A2(n126), .B1(B[7]), .B2(n128), .ZN(n37) );
  INV_X1 U70 ( .A(n36), .ZN(Y[8]) );
  AOI22_X1 U71 ( .A1(A[8]), .A2(n126), .B1(B[8]), .B2(n128), .ZN(n36) );
  INV_X1 U72 ( .A(n34), .ZN(Y[9]) );
  AOI22_X1 U73 ( .A1(A[9]), .A2(n127), .B1(n135), .B2(B[9]), .ZN(n34) );
  INV_X1 U74 ( .A(n42), .ZN(Y[31]) );
  AOI22_X1 U75 ( .A1(A[31]), .A2(n127), .B1(B[31]), .B2(n129), .ZN(n42) );
  BUF_X1 U76 ( .A(SEL), .Z(n125) );
  BUF_X1 U77 ( .A(SEL), .Z(n124) );
  BUF_X1 U78 ( .A(SEL), .Z(n123) );
endmodule


module registro_N32_3 ( data, enable, clock, clear, Q );
  input [31:0] data;
  output [31:0] Q;
  input enable, clock, clear;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net44624, net44625, net44626, net44627, net44628, net44629,
         net44630, net44631, net44632, net44633, net44634, net44635, net44636,
         net44637, net44638, net44639, net44640, net44641, net44642, net44643,
         net44644, net44645, net44646, net44647, net44648, net44649, net44650,
         net44651, net44652, net44653, net103958, net103959, net120727, n132,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148;
  assign Q[30] = net103958;
  assign Q[31] = net103959;
  assign n132 = clear;

  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(clock), .RN(n140), .Q(Q[27]), .QN(net44651) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(clock), .RN(n140), .Q(Q[26]), .QN(net44650) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(clock), .RN(n141), .Q(Q[25]), .QN(net44649) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(clock), .RN(n141), .Q(Q[24]), .QN(net44648) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(clock), .RN(n141), .Q(Q[23]), .QN(net44647) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(clock), .RN(n141), .Q(Q[22]), .QN(
        net44646) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(clock), .RN(n140), .Q(Q[21]), .QN(
        net44645) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(clock), .RN(n142), .Q(Q[20]), .QN(
        net44644) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(clock), .RN(n140), .Q(Q[19]), .QN(
        net44643) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(clock), .RN(n141), .Q(Q[18]), .QN(
        net44642) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(clock), .RN(n141), .Q(Q[17]), .QN(
        net44641) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(clock), .RN(n141), .Q(Q[16]), .QN(
        net44640) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(clock), .RN(n140), .Q(Q[15]), .QN(
        net44639) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(clock), .RN(n140), .Q(Q[14]), .QN(
        net44638) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(clock), .RN(n141), .Q(Q[13]), .QN(
        net44637) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(clock), .RN(n140), .Q(Q[12]), .QN(
        net44636) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(clock), .RN(n140), .Q(Q[11]), .QN(
        net44635) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(clock), .RN(n141), .Q(Q[10]), .QN(
        net44634) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(clock), .RN(n141), .Q(Q[9]), .QN(net44633)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(clock), .RN(n142), .Q(Q[8]), .QN(net44632)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(clock), .RN(n141), .Q(Q[7]), .QN(net44631)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(clock), .RN(n140), .Q(Q[6]), .QN(net44630)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(clock), .RN(n141), .Q(Q[5]), .QN(net44629)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(clock), .RN(n140), .Q(Q[4]), .QN(net44628)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(clock), .RN(n142), .Q(Q[3]), .QN(net44627)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(clock), .RN(n142), .Q(Q[2]), .QN(net44626)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(clock), .RN(n140), .Q(Q[1]), .QN(net44625)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(clock), .RN(n140), .Q(Q[0]), .QN(net44624)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(clock), .RN(n141), .Q(Q[29]), .QN(net44653) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(clock), .RN(n141), .Q(net103958), .QN(
        net120727) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(clock), .RN(n140), .Q(Q[28]), .QN(net44652) );
  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(clock), .RN(n140), .Q(net103959) );
  INV_X1 U2 ( .A(enable), .ZN(n139) );
  MUX2_X1 U3 ( .A(data[31]), .B(net103959), .S(n139), .Z(n1) );
  BUF_X1 U4 ( .A(n132), .Z(n141) );
  BUF_X1 U5 ( .A(n132), .Z(n140) );
  BUF_X1 U6 ( .A(n132), .Z(n142) );
  OAI21_X1 U7 ( .B1(net44642), .B2(n147), .A(n59), .ZN(n14) );
  NAND2_X1 U8 ( .A1(data[18]), .A2(n143), .ZN(n59) );
  OAI21_X1 U9 ( .B1(net44648), .B2(n145), .A(n34), .ZN(n8) );
  NAND2_X1 U10 ( .A1(data[24]), .A2(n143), .ZN(n34) );
  OAI21_X1 U11 ( .B1(net44649), .B2(n145), .A(n35), .ZN(n7) );
  NAND2_X1 U12 ( .A1(data[25]), .A2(n143), .ZN(n35) );
  OAI21_X1 U13 ( .B1(net44653), .B2(n146), .A(n42), .ZN(n3) );
  NAND2_X1 U14 ( .A1(data[29]), .A2(n145), .ZN(n42) );
  OAI21_X1 U15 ( .B1(net44643), .B2(n147), .A(n60), .ZN(n13) );
  NAND2_X1 U16 ( .A1(data[19]), .A2(n143), .ZN(n60) );
  OAI21_X1 U17 ( .B1(net44636), .B2(n147), .A(n52), .ZN(n20) );
  NAND2_X1 U18 ( .A1(data[12]), .A2(n144), .ZN(n52) );
  OAI21_X1 U19 ( .B1(net44645), .B2(n148), .A(n62), .ZN(n11) );
  NAND2_X1 U20 ( .A1(data[21]), .A2(n143), .ZN(n62) );
  OAI21_X1 U21 ( .B1(net44639), .B2(n147), .A(n56), .ZN(n17) );
  NAND2_X1 U22 ( .A1(data[15]), .A2(n144), .ZN(n56) );
  OAI21_X1 U23 ( .B1(net44652), .B2(n145), .A(n38), .ZN(n4) );
  NAND2_X1 U24 ( .A1(data[28]), .A2(n144), .ZN(n38) );
  OAI21_X1 U25 ( .B1(net44651), .B2(n145), .A(n37), .ZN(n5) );
  NAND2_X1 U26 ( .A1(data[27]), .A2(n143), .ZN(n37) );
  OAI21_X1 U27 ( .B1(net120727), .B2(n147), .A(n53), .ZN(n2) );
  NAND2_X1 U28 ( .A1(data[30]), .A2(n144), .ZN(n53) );
  OAI21_X1 U29 ( .B1(net44650), .B2(n146), .A(n36), .ZN(n6) );
  NAND2_X1 U30 ( .A1(data[26]), .A2(n143), .ZN(n36) );
  OAI21_X1 U31 ( .B1(net44647), .B2(n146), .A(n33), .ZN(n9) );
  NAND2_X1 U32 ( .A1(n148), .A2(data[23]), .ZN(n33) );
  OAI21_X1 U33 ( .B1(net44646), .B2(n148), .A(n63), .ZN(n10) );
  NAND2_X1 U34 ( .A1(data[22]), .A2(n143), .ZN(n63) );
  OAI21_X1 U35 ( .B1(net44644), .B2(n148), .A(n61), .ZN(n12) );
  NAND2_X1 U36 ( .A1(data[20]), .A2(n143), .ZN(n61) );
  OAI21_X1 U37 ( .B1(net44638), .B2(n147), .A(n55), .ZN(n18) );
  NAND2_X1 U38 ( .A1(data[14]), .A2(n144), .ZN(n55) );
  OAI21_X1 U39 ( .B1(net44641), .B2(n147), .A(n58), .ZN(n15) );
  NAND2_X1 U40 ( .A1(data[17]), .A2(n143), .ZN(n58) );
  OAI21_X1 U41 ( .B1(net44637), .B2(n147), .A(n54), .ZN(n19) );
  NAND2_X1 U42 ( .A1(data[13]), .A2(n144), .ZN(n54) );
  OAI21_X1 U43 ( .B1(net44640), .B2(n147), .A(n57), .ZN(n16) );
  NAND2_X1 U44 ( .A1(data[16]), .A2(n143), .ZN(n57) );
  OAI21_X1 U45 ( .B1(net44629), .B2(n146), .A(n45), .ZN(n27) );
  NAND2_X1 U46 ( .A1(data[5]), .A2(n145), .ZN(n45) );
  OAI21_X1 U47 ( .B1(net44632), .B2(n146), .A(n48), .ZN(n24) );
  NAND2_X1 U48 ( .A1(data[8]), .A2(n145), .ZN(n48) );
  OAI21_X1 U49 ( .B1(net44630), .B2(n146), .A(n46), .ZN(n26) );
  NAND2_X1 U50 ( .A1(data[6]), .A2(n145), .ZN(n46) );
  OAI21_X1 U51 ( .B1(net44635), .B2(n147), .A(n51), .ZN(n21) );
  NAND2_X1 U52 ( .A1(data[11]), .A2(n144), .ZN(n51) );
  OAI21_X1 U53 ( .B1(net44631), .B2(n146), .A(n47), .ZN(n25) );
  NAND2_X1 U54 ( .A1(data[7]), .A2(n145), .ZN(n47) );
  OAI21_X1 U55 ( .B1(net44633), .B2(n147), .A(n49), .ZN(n23) );
  NAND2_X1 U56 ( .A1(data[9]), .A2(n145), .ZN(n49) );
  OAI21_X1 U57 ( .B1(net44634), .B2(n147), .A(n50), .ZN(n22) );
  NAND2_X1 U58 ( .A1(data[10]), .A2(n144), .ZN(n50) );
  OAI21_X1 U59 ( .B1(net44627), .B2(n146), .A(n43), .ZN(n29) );
  NAND2_X1 U60 ( .A1(data[3]), .A2(n144), .ZN(n43) );
  OAI21_X1 U61 ( .B1(net44626), .B2(n146), .A(n41), .ZN(n30) );
  NAND2_X1 U62 ( .A1(data[2]), .A2(n144), .ZN(n41) );
  OAI21_X1 U63 ( .B1(net44624), .B2(n146), .A(n39), .ZN(n32) );
  NAND2_X1 U64 ( .A1(data[0]), .A2(n144), .ZN(n39) );
  OAI21_X1 U65 ( .B1(net44625), .B2(n145), .A(n40), .ZN(n31) );
  NAND2_X1 U66 ( .A1(data[1]), .A2(n144), .ZN(n40) );
  OAI21_X1 U67 ( .B1(net44628), .B2(n146), .A(n44), .ZN(n28) );
  NAND2_X1 U68 ( .A1(data[4]), .A2(n145), .ZN(n44) );
  CLKBUF_X1 U69 ( .A(enable), .Z(n143) );
  CLKBUF_X1 U70 ( .A(enable), .Z(n144) );
  CLKBUF_X1 U71 ( .A(enable), .Z(n145) );
  CLKBUF_X1 U72 ( .A(enable), .Z(n146) );
  CLKBUF_X1 U73 ( .A(enable), .Z(n147) );
  CLKBUF_X1 U74 ( .A(enable), .Z(n148) );
endmodule


module registro_N5_2 ( data, enable, clock, clear, Q );
  input [4:0] data;
  output [4:0] Q;
  input enable, clock, clear;
  wire   n1, n2, n3, n4, n5, net44880, net44881, net44882, net44883, net44884,
         n6, n7, n8, n9, n10;

  DFFR_X1 \Q_reg[4]  ( .D(n1), .CK(clock), .RN(clear), .Q(Q[4]), .QN(net44884)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n2), .CK(clock), .RN(clear), .Q(Q[3]), .QN(net44883)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n3), .CK(clock), .RN(clear), .Q(Q[2]), .QN(net44882)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n4), .CK(clock), .RN(clear), .Q(Q[1]), .QN(net44881)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n5), .CK(clock), .RN(clear), .Q(Q[0]), .QN(net44880)
         );
  OAI21_X1 U2 ( .B1(net44880), .B2(enable), .A(n6), .ZN(n5) );
  NAND2_X1 U3 ( .A1(enable), .A2(data[0]), .ZN(n6) );
  OAI21_X1 U4 ( .B1(net44881), .B2(enable), .A(n7), .ZN(n4) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(enable), .ZN(n7) );
  OAI21_X1 U6 ( .B1(net44882), .B2(enable), .A(n8), .ZN(n3) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(enable), .ZN(n8) );
  OAI21_X1 U8 ( .B1(net44883), .B2(enable), .A(n9), .ZN(n2) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(enable), .ZN(n9) );
  OAI21_X1 U10 ( .B1(net44884), .B2(enable), .A(n10), .ZN(n1) );
  NAND2_X1 U11 ( .A1(data[4]), .A2(enable), .ZN(n10) );
endmodule


module registro_N32_4 ( data, enable, clock, clear, Q );
  input [31:0] data;
  output [31:0] Q;
  input enable, clock, clear;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net44624, net44625, net44626, net44627, net44628, net44629,
         net44630, net44631, net44632, net44633, net44634, net44635, net44636,
         net44637, net44638, net44639, net44640, net44641, net44642, net44643,
         net44644, net44645, net44646, net44647, net44648, net44649, net44650,
         net44651, net44652, net44653, net44654, net44655, n135, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n142, n143, n144, n145, n146, n147, n148, n149, n150;
  assign n135 = clear;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(clock), .RN(n144), .Q(Q[31]), .QN(net44655) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(clock), .RN(n144), .Q(Q[30]), .QN(net44654) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(clock), .RN(n144), .Q(Q[29]), .QN(net44653) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(clock), .RN(n144), .Q(Q[28]), .QN(net44652) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(clock), .RN(n144), .Q(Q[27]), .QN(net44651) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(clock), .RN(n144), .Q(Q[26]), .QN(net44650) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(clock), .RN(n144), .Q(Q[25]), .QN(net44649) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(clock), .RN(n144), .Q(Q[24]), .QN(net44648) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(clock), .RN(n144), .Q(Q[23]), .QN(net44647) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(clock), .RN(n144), .Q(Q[22]), .QN(
        net44646) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(clock), .RN(n142), .Q(Q[21]), .QN(
        net44645) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(clock), .RN(n142), .Q(Q[20]), .QN(
        net44644) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(clock), .RN(n142), .Q(Q[19]), .QN(
        net44643) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(clock), .RN(n142), .Q(Q[18]), .QN(
        net44642) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(clock), .RN(n142), .Q(Q[17]), .QN(
        net44641) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(clock), .RN(n142), .Q(Q[16]), .QN(
        net44640) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(clock), .RN(n142), .Q(Q[15]), .QN(
        net44639) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(clock), .RN(n142), .Q(Q[14]), .QN(
        net44638) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(clock), .RN(n142), .Q(Q[13]), .QN(
        net44637) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(clock), .RN(n142), .Q(Q[12]), .QN(
        net44636) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(clock), .RN(n142), .Q(Q[11]), .QN(
        net44635) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(clock), .RN(n143), .Q(Q[10]), .QN(
        net44634) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(clock), .RN(n143), .Q(Q[9]), .QN(net44633)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(clock), .RN(n143), .Q(Q[8]), .QN(net44632)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(clock), .RN(n143), .Q(Q[7]), .QN(net44631)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(clock), .RN(n143), .Q(Q[6]), .QN(net44630)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(clock), .RN(n143), .Q(Q[5]), .QN(net44629)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(clock), .RN(n143), .Q(Q[4]), .QN(net44628)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(clock), .RN(n143), .Q(Q[3]), .QN(net44627)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(clock), .RN(n143), .Q(Q[2]), .QN(net44626)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(clock), .RN(n143), .Q(Q[1]), .QN(net44625)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(clock), .RN(n143), .Q(Q[0]), .QN(net44624)
         );
  BUF_X1 U2 ( .A(n135), .Z(n143) );
  BUF_X1 U3 ( .A(n135), .Z(n142) );
  BUF_X1 U4 ( .A(n135), .Z(n144) );
  BUF_X1 U5 ( .A(enable), .Z(n146) );
  BUF_X1 U6 ( .A(enable), .Z(n145) );
  BUF_X1 U7 ( .A(enable), .Z(n147) );
  BUF_X1 U8 ( .A(enable), .Z(n149) );
  BUF_X1 U9 ( .A(enable), .Z(n148) );
  OAI21_X1 U10 ( .B1(net44625), .B2(n147), .A(n40), .ZN(n31) );
  NAND2_X1 U11 ( .A1(data[1]), .A2(n146), .ZN(n40) );
  OAI21_X1 U12 ( .B1(net44648), .B2(n147), .A(n34), .ZN(n8) );
  NAND2_X1 U13 ( .A1(data[24]), .A2(n145), .ZN(n34) );
  OAI21_X1 U14 ( .B1(net44649), .B2(n147), .A(n35), .ZN(n7) );
  NAND2_X1 U15 ( .A1(data[25]), .A2(n145), .ZN(n35) );
  OAI21_X1 U16 ( .B1(net44651), .B2(n147), .A(n37), .ZN(n5) );
  NAND2_X1 U17 ( .A1(data[27]), .A2(n145), .ZN(n37) );
  OAI21_X1 U18 ( .B1(net44652), .B2(n147), .A(n38), .ZN(n4) );
  NAND2_X1 U19 ( .A1(data[28]), .A2(n146), .ZN(n38) );
  OAI21_X1 U20 ( .B1(net44624), .B2(n148), .A(n39), .ZN(n32) );
  NAND2_X1 U21 ( .A1(data[0]), .A2(n146), .ZN(n39) );
  OAI21_X1 U22 ( .B1(net44626), .B2(n148), .A(n41), .ZN(n30) );
  NAND2_X1 U23 ( .A1(data[2]), .A2(n146), .ZN(n41) );
  OAI21_X1 U24 ( .B1(net44627), .B2(n148), .A(n43), .ZN(n29) );
  NAND2_X1 U25 ( .A1(data[3]), .A2(n146), .ZN(n43) );
  OAI21_X1 U26 ( .B1(net44634), .B2(n149), .A(n50), .ZN(n22) );
  NAND2_X1 U27 ( .A1(data[10]), .A2(n146), .ZN(n50) );
  OAI21_X1 U28 ( .B1(net44635), .B2(n149), .A(n51), .ZN(n21) );
  NAND2_X1 U29 ( .A1(data[11]), .A2(n146), .ZN(n51) );
  OAI21_X1 U30 ( .B1(net44636), .B2(n149), .A(n52), .ZN(n20) );
  NAND2_X1 U31 ( .A1(data[12]), .A2(n146), .ZN(n52) );
  OAI21_X1 U32 ( .B1(net44637), .B2(n149), .A(n54), .ZN(n19) );
  NAND2_X1 U33 ( .A1(data[13]), .A2(n146), .ZN(n54) );
  OAI21_X1 U34 ( .B1(net44638), .B2(n149), .A(n55), .ZN(n18) );
  NAND2_X1 U35 ( .A1(data[14]), .A2(n146), .ZN(n55) );
  OAI21_X1 U36 ( .B1(net44639), .B2(n149), .A(n56), .ZN(n17) );
  NAND2_X1 U37 ( .A1(data[15]), .A2(n146), .ZN(n56) );
  OAI21_X1 U38 ( .B1(net44640), .B2(n149), .A(n57), .ZN(n16) );
  NAND2_X1 U39 ( .A1(data[16]), .A2(n145), .ZN(n57) );
  OAI21_X1 U40 ( .B1(net44641), .B2(n149), .A(n58), .ZN(n15) );
  NAND2_X1 U41 ( .A1(data[17]), .A2(n145), .ZN(n58) );
  OAI21_X1 U42 ( .B1(net44642), .B2(n149), .A(n59), .ZN(n14) );
  NAND2_X1 U43 ( .A1(data[18]), .A2(n145), .ZN(n59) );
  OAI21_X1 U44 ( .B1(net44643), .B2(n149), .A(n60), .ZN(n13) );
  NAND2_X1 U45 ( .A1(data[19]), .A2(n145), .ZN(n60) );
  OAI21_X1 U46 ( .B1(net44647), .B2(n148), .A(n33), .ZN(n9) );
  NAND2_X1 U47 ( .A1(n150), .A2(data[23]), .ZN(n33) );
  OAI21_X1 U48 ( .B1(net44650), .B2(n148), .A(n36), .ZN(n6) );
  NAND2_X1 U49 ( .A1(data[26]), .A2(n145), .ZN(n36) );
  OAI21_X1 U50 ( .B1(net44654), .B2(n149), .A(n53), .ZN(n2) );
  NAND2_X1 U51 ( .A1(data[30]), .A2(n146), .ZN(n53) );
  OAI21_X1 U52 ( .B1(net44655), .B2(n148), .A(n64), .ZN(n1) );
  NAND2_X1 U53 ( .A1(data[31]), .A2(n145), .ZN(n64) );
  OAI21_X1 U54 ( .B1(net44644), .B2(n150), .A(n61), .ZN(n12) );
  NAND2_X1 U55 ( .A1(data[20]), .A2(n145), .ZN(n61) );
  OAI21_X1 U56 ( .B1(net44645), .B2(n150), .A(n62), .ZN(n11) );
  NAND2_X1 U57 ( .A1(data[21]), .A2(n145), .ZN(n62) );
  OAI21_X1 U58 ( .B1(net44646), .B2(n150), .A(n63), .ZN(n10) );
  NAND2_X1 U59 ( .A1(data[22]), .A2(n145), .ZN(n63) );
  OAI21_X1 U60 ( .B1(net44628), .B2(n148), .A(n44), .ZN(n28) );
  NAND2_X1 U61 ( .A1(data[4]), .A2(n147), .ZN(n44) );
  OAI21_X1 U62 ( .B1(net44629), .B2(n148), .A(n45), .ZN(n27) );
  NAND2_X1 U63 ( .A1(data[5]), .A2(n147), .ZN(n45) );
  OAI21_X1 U64 ( .B1(net44630), .B2(n148), .A(n46), .ZN(n26) );
  NAND2_X1 U65 ( .A1(data[6]), .A2(n147), .ZN(n46) );
  OAI21_X1 U66 ( .B1(net44631), .B2(n148), .A(n47), .ZN(n25) );
  NAND2_X1 U67 ( .A1(data[7]), .A2(n147), .ZN(n47) );
  OAI21_X1 U68 ( .B1(net44632), .B2(n148), .A(n48), .ZN(n24) );
  NAND2_X1 U69 ( .A1(data[8]), .A2(n147), .ZN(n48) );
  OAI21_X1 U70 ( .B1(net44633), .B2(n149), .A(n49), .ZN(n23) );
  NAND2_X1 U71 ( .A1(data[9]), .A2(n147), .ZN(n49) );
  OAI21_X1 U72 ( .B1(net44653), .B2(n148), .A(n42), .ZN(n3) );
  NAND2_X1 U73 ( .A1(data[29]), .A2(n147), .ZN(n42) );
  CLKBUF_X1 U74 ( .A(enable), .Z(n150) );
endmodule


module registro_N32_5 ( data, enable, clock, clear, Q );
  input [31:0] data;
  output [31:0] Q;
  input enable, clock, clear;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net44624, net44625, net44626, net44627, net44628, net44629,
         net44630, net44631, net44632, net44633, net44634, net44635, net44636,
         net44637, net44638, net44639, net44640, net44641, net44642, net44643,
         net44644, net44645, net44646, net44647, net44648, net44649, net44650,
         net44651, net44652, net44653, net44654, net44655, n136, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n143, n144, n145, n146, n147, n148, n149, n150, n151;
  assign n136 = clear;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(clock), .RN(n145), .Q(Q[31]), .QN(net44655) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(clock), .RN(n145), .Q(Q[30]), .QN(net44654) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(clock), .RN(n145), .Q(Q[29]), .QN(net44653) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(clock), .RN(n145), .Q(Q[28]), .QN(net44652) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(clock), .RN(n145), .Q(Q[27]), .QN(net44651) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(clock), .RN(n145), .Q(Q[26]), .QN(net44650) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(clock), .RN(n145), .Q(Q[25]), .QN(net44649) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(clock), .RN(n145), .Q(Q[24]), .QN(net44648) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(clock), .RN(n145), .Q(Q[23]), .QN(net44647) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(clock), .RN(n145), .Q(Q[22]), .QN(
        net44646) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(clock), .RN(n143), .Q(Q[21]), .QN(
        net44645) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(clock), .RN(n143), .Q(Q[20]), .QN(
        net44644) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(clock), .RN(n143), .Q(Q[19]), .QN(
        net44643) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(clock), .RN(n143), .Q(Q[18]), .QN(
        net44642) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(clock), .RN(n143), .Q(Q[17]), .QN(
        net44641) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(clock), .RN(n143), .Q(Q[16]), .QN(
        net44640) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(clock), .RN(n143), .Q(Q[15]), .QN(
        net44639) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(clock), .RN(n143), .Q(Q[14]), .QN(
        net44638) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(clock), .RN(n143), .Q(Q[13]), .QN(
        net44637) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(clock), .RN(n143), .Q(Q[12]), .QN(
        net44636) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(clock), .RN(n143), .Q(Q[11]), .QN(
        net44635) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(clock), .RN(n144), .Q(Q[10]), .QN(
        net44634) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(clock), .RN(n144), .Q(Q[9]), .QN(net44633)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(clock), .RN(n144), .Q(Q[8]), .QN(net44632)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(clock), .RN(n144), .Q(Q[7]), .QN(net44631)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(clock), .RN(n144), .Q(Q[6]), .QN(net44630)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(clock), .RN(n144), .Q(Q[5]), .QN(net44629)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(clock), .RN(n144), .Q(Q[4]), .QN(net44628)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(clock), .RN(n144), .Q(Q[3]), .QN(net44627)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(clock), .RN(n144), .Q(Q[2]), .QN(net44626)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(clock), .RN(n144), .Q(Q[1]), .QN(net44625)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(clock), .RN(n144), .Q(Q[0]), .QN(net44624)
         );
  CLKBUF_X1 U2 ( .A(enable), .Z(n149) );
  BUF_X1 U3 ( .A(n136), .Z(n144) );
  BUF_X1 U4 ( .A(n136), .Z(n143) );
  BUF_X1 U5 ( .A(n136), .Z(n145) );
  OAI21_X1 U6 ( .B1(net44625), .B2(n148), .A(n40), .ZN(n31) );
  NAND2_X1 U7 ( .A1(data[1]), .A2(n147), .ZN(n40) );
  OAI21_X1 U8 ( .B1(net44648), .B2(n148), .A(n34), .ZN(n8) );
  NAND2_X1 U9 ( .A1(data[24]), .A2(n146), .ZN(n34) );
  OAI21_X1 U10 ( .B1(net44649), .B2(n148), .A(n35), .ZN(n7) );
  NAND2_X1 U11 ( .A1(data[25]), .A2(n146), .ZN(n35) );
  OAI21_X1 U12 ( .B1(net44651), .B2(n148), .A(n37), .ZN(n5) );
  NAND2_X1 U13 ( .A1(data[27]), .A2(n146), .ZN(n37) );
  OAI21_X1 U14 ( .B1(net44652), .B2(n148), .A(n38), .ZN(n4) );
  NAND2_X1 U15 ( .A1(data[28]), .A2(n147), .ZN(n38) );
  OAI21_X1 U16 ( .B1(net44626), .B2(n149), .A(n41), .ZN(n30) );
  NAND2_X1 U17 ( .A1(data[2]), .A2(n147), .ZN(n41) );
  OAI21_X1 U18 ( .B1(net44629), .B2(n149), .A(n45), .ZN(n27) );
  NAND2_X1 U19 ( .A1(data[5]), .A2(n148), .ZN(n45) );
  OAI21_X1 U20 ( .B1(net44654), .B2(n150), .A(n53), .ZN(n2) );
  NAND2_X1 U21 ( .A1(data[30]), .A2(n147), .ZN(n53) );
  OAI21_X1 U22 ( .B1(net44630), .B2(n149), .A(n46), .ZN(n26) );
  NAND2_X1 U23 ( .A1(data[6]), .A2(n148), .ZN(n46) );
  OAI21_X1 U24 ( .B1(net44631), .B2(n149), .A(n47), .ZN(n25) );
  NAND2_X1 U25 ( .A1(data[7]), .A2(n148), .ZN(n47) );
  OAI21_X1 U26 ( .B1(net44628), .B2(n149), .A(n44), .ZN(n28) );
  NAND2_X1 U27 ( .A1(data[4]), .A2(n148), .ZN(n44) );
  OAI21_X1 U28 ( .B1(net44655), .B2(n149), .A(n64), .ZN(n1) );
  NAND2_X1 U29 ( .A1(data[31]), .A2(n146), .ZN(n64) );
  OAI21_X1 U30 ( .B1(net44627), .B2(n149), .A(n43), .ZN(n29) );
  NAND2_X1 U31 ( .A1(data[3]), .A2(n147), .ZN(n43) );
  OAI21_X1 U32 ( .B1(net44647), .B2(n149), .A(n33), .ZN(n9) );
  NAND2_X1 U33 ( .A1(n151), .A2(data[23]), .ZN(n33) );
  OAI21_X1 U34 ( .B1(net44624), .B2(n149), .A(n39), .ZN(n32) );
  NAND2_X1 U35 ( .A1(data[0]), .A2(n147), .ZN(n39) );
  OAI21_X1 U36 ( .B1(net44634), .B2(n150), .A(n50), .ZN(n22) );
  NAND2_X1 U37 ( .A1(data[10]), .A2(n147), .ZN(n50) );
  OAI21_X1 U38 ( .B1(net44635), .B2(n150), .A(n51), .ZN(n21) );
  NAND2_X1 U39 ( .A1(data[11]), .A2(n147), .ZN(n51) );
  OAI21_X1 U40 ( .B1(net44636), .B2(n150), .A(n52), .ZN(n20) );
  NAND2_X1 U41 ( .A1(data[12]), .A2(n147), .ZN(n52) );
  OAI21_X1 U42 ( .B1(net44637), .B2(n150), .A(n54), .ZN(n19) );
  NAND2_X1 U43 ( .A1(data[13]), .A2(n147), .ZN(n54) );
  OAI21_X1 U44 ( .B1(net44638), .B2(n150), .A(n55), .ZN(n18) );
  NAND2_X1 U45 ( .A1(data[14]), .A2(n147), .ZN(n55) );
  OAI21_X1 U46 ( .B1(net44639), .B2(n150), .A(n56), .ZN(n17) );
  NAND2_X1 U47 ( .A1(data[15]), .A2(n147), .ZN(n56) );
  OAI21_X1 U48 ( .B1(net44640), .B2(n150), .A(n57), .ZN(n16) );
  NAND2_X1 U49 ( .A1(data[16]), .A2(n146), .ZN(n57) );
  OAI21_X1 U50 ( .B1(net44641), .B2(n150), .A(n58), .ZN(n15) );
  NAND2_X1 U51 ( .A1(data[17]), .A2(n146), .ZN(n58) );
  OAI21_X1 U52 ( .B1(net44642), .B2(n150), .A(n59), .ZN(n14) );
  NAND2_X1 U53 ( .A1(data[18]), .A2(n146), .ZN(n59) );
  OAI21_X1 U54 ( .B1(net44643), .B2(n150), .A(n60), .ZN(n13) );
  NAND2_X1 U55 ( .A1(data[19]), .A2(n146), .ZN(n60) );
  OAI21_X1 U56 ( .B1(net44650), .B2(n149), .A(n36), .ZN(n6) );
  NAND2_X1 U57 ( .A1(data[26]), .A2(n146), .ZN(n36) );
  OAI21_X1 U58 ( .B1(net44632), .B2(n149), .A(n48), .ZN(n24) );
  NAND2_X1 U59 ( .A1(data[8]), .A2(n148), .ZN(n48) );
  OAI21_X1 U60 ( .B1(net44633), .B2(n150), .A(n49), .ZN(n23) );
  NAND2_X1 U61 ( .A1(data[9]), .A2(n148), .ZN(n49) );
  OAI21_X1 U62 ( .B1(net44653), .B2(n149), .A(n42), .ZN(n3) );
  NAND2_X1 U63 ( .A1(data[29]), .A2(n148), .ZN(n42) );
  OAI21_X1 U64 ( .B1(net44644), .B2(n151), .A(n61), .ZN(n12) );
  NAND2_X1 U65 ( .A1(data[20]), .A2(n146), .ZN(n61) );
  OAI21_X1 U66 ( .B1(net44645), .B2(n151), .A(n62), .ZN(n11) );
  NAND2_X1 U67 ( .A1(data[21]), .A2(n146), .ZN(n62) );
  OAI21_X1 U68 ( .B1(net44646), .B2(n151), .A(n63), .ZN(n10) );
  NAND2_X1 U69 ( .A1(data[22]), .A2(n146), .ZN(n63) );
  BUF_X1 U70 ( .A(enable), .Z(n147) );
  BUF_X1 U71 ( .A(enable), .Z(n146) );
  BUF_X1 U72 ( .A(enable), .Z(n148) );
  BUF_X1 U73 ( .A(enable), .Z(n150) );
  CLKBUF_X1 U74 ( .A(enable), .Z(n151) );
endmodule


module AluOpCodeGen ( IR_opcode, IR_func, AluOpCode, Add_Subn, CompareCode, 
        ShiftOpCode );
  input [5:0] IR_opcode;
  input [10:0] IR_func;
  output [2:0] AluOpCode;
  output [3:0] CompareCode;
  output [2:0] ShiftOpCode;
  output Add_Subn;
  wire   n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43;
  assign ShiftOpCode[2] = ShiftOpCode[0];

  OAI33_X1 U40 ( .A1(n27), .A2(n17), .A3(n35), .B1(n31), .B2(n20), .B3(n36), 
        .ZN(n34) );
  NAND3_X1 U41 ( .A1(n26), .A2(n29), .A3(IR_func[2]), .ZN(n37) );
  OAI33_X1 U42 ( .A1(n27), .A2(IR_func[2]), .A3(n35), .B1(n31), .B2(
        IR_opcode[2]), .B3(n36), .ZN(Add_Subn) );
  NAND3_X1 U43 ( .A1(n39), .A2(n32), .A3(n16), .ZN(n40) );
  INV_X1 U3 ( .A(ShiftOpCode[0]), .ZN(n25) );
  OAI21_X1 U4 ( .B1(n17), .B2(n18), .A(n19), .ZN(CompareCode[1]) );
  OAI221_X1 U5 ( .B1(n20), .B2(n36), .C1(n17), .C2(n35), .A(n25), .ZN(
        AluOpCode[0]) );
  OAI211_X1 U6 ( .C1(n24), .C2(n22), .A(n18), .B(n25), .ZN(AluOpCode[2]) );
  NOR3_X1 U7 ( .A1(n16), .A2(n15), .A3(n39), .ZN(n21) );
  NAND2_X1 U8 ( .A1(n13), .A2(n14), .ZN(ShiftOpCode[0]) );
  OR3_X1 U9 ( .A1(n20), .A2(n40), .A3(n24), .ZN(n13) );
  OR3_X1 U10 ( .A1(n20), .A2(n21), .A3(n22), .ZN(n19) );
  NOR3_X1 U11 ( .A1(n15), .A2(IR_opcode[3]), .A3(IR_opcode[0]), .ZN(
        CompareCode[3]) );
  NOR4_X1 U12 ( .A1(IR_func[10]), .A2(n40), .A3(n41), .A4(n42), .ZN(n26) );
  OR3_X1 U13 ( .A1(IR_func[7]), .A2(IR_func[6]), .A3(IR_func[4]), .ZN(n41) );
  NAND4_X1 U14 ( .A1(n20), .A2(n24), .A3(n31), .A4(n43), .ZN(n42) );
  NOR2_X1 U15 ( .A1(IR_func[9]), .A2(IR_func[8]), .ZN(n43) );
  NAND4_X1 U16 ( .A1(IR_func[5]), .A2(n26), .A3(n38), .A4(n29), .ZN(n35) );
  INV_X1 U17 ( .A(IR_opcode[4]), .ZN(n24) );
  INV_X1 U18 ( .A(IR_opcode[2]), .ZN(n20) );
  INV_X1 U19 ( .A(IR_opcode[1]), .ZN(n31) );
  INV_X1 U20 ( .A(IR_opcode[5]), .ZN(n32) );
  INV_X1 U21 ( .A(IR_opcode[0]), .ZN(n16) );
  INV_X1 U22 ( .A(IR_opcode[3]), .ZN(n39) );
  OAI22_X1 U23 ( .A1(IR_opcode[1]), .A2(n13), .B1(IR_func[1]), .B2(n14), .ZN(
        ShiftOpCode[1]) );
  NAND4_X1 U24 ( .A1(n26), .A2(n27), .A3(IR_func[0]), .A4(n28), .ZN(n18) );
  NOR2_X1 U25 ( .A1(n29), .A2(n30), .ZN(n28) );
  NAND4_X1 U26 ( .A1(IR_opcode[3]), .A2(IR_opcode[0]), .A3(n31), .A4(n32), 
        .ZN(n22) );
  NAND4_X1 U27 ( .A1(IR_opcode[2]), .A2(n31), .A3(n24), .A4(n32), .ZN(n15) );
  NOR3_X1 U28 ( .A1(n16), .A2(IR_opcode[3]), .A3(n15), .ZN(CompareCode[2]) );
  NAND4_X1 U29 ( .A1(IR_opcode[3]), .A2(n16), .A3(n24), .A4(n32), .ZN(n36) );
  OAI21_X1 U30 ( .B1(IR_func[2]), .B2(n18), .A(n23), .ZN(CompareCode[0]) );
  OR3_X1 U31 ( .A1(n24), .A2(IR_opcode[2]), .A3(n22), .ZN(n23) );
  OR3_X1 U32 ( .A1(n21), .A2(n33), .A3(n34), .ZN(AluOpCode[1]) );
  NOR4_X1 U33 ( .A1(IR_func[1]), .A2(n37), .A3(n38), .A4(n30), .ZN(n33) );
  INV_X1 U34 ( .A(IR_func[3]), .ZN(n29) );
  INV_X1 U35 ( .A(IR_func[2]), .ZN(n17) );
  OR3_X1 U36 ( .A1(IR_func[0]), .A2(IR_func[5]), .A3(n37), .ZN(n14) );
  INV_X1 U37 ( .A(IR_func[1]), .ZN(n27) );
  INV_X1 U38 ( .A(IR_func[0]), .ZN(n38) );
  INV_X1 U39 ( .A(IR_func[5]), .ZN(n30) );
endmodule


module ALU_N32 ( AluOpCode, CompareOpCode, Add_subn, ShiftOpCode, DATA1, DATA2, 
        OUTALU, return_address, CompBranch );
  input [2:0] AluOpCode;
  input [3:0] CompareOpCode;
  input [2:0] ShiftOpCode;
  input [31:0] DATA1;
  input [31:0] DATA2;
  output [31:0] OUTALU;
  output [31:0] return_address;
  input Add_subn;
  output CompBranch;
  wire   comp_eq, comp_greater, sel_mux_comp_out, n58, n71, n72, n74, n89, n91,
         n100, n102, n111, n123, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n3, n4, n5, n146, n147, n148, n149, n150, n151, n152,
         n153, n154, n155, n156, n157, n158, n159, n160, n161, n162, n163,
         n164, n165, n166, n167, n168, n169, n170, n171;
  wire   [31:0] shift_out;
  wire   [31:0] AND_OUT;
  wire   [31:0] OR_OUT;
  wire   [31:0] XOR_OUT;
  wire   [31:0] add_sub_out;
  wire   [31:0] comp_out;
  assign n58 = DATA2[0];
  assign n71 = DATA1[6];
  assign n72 = DATA1[7];
  assign n74 = DATA1[9];
  assign n89 = DATA1[27];
  assign n91 = DATA1[30];
  assign n100 = DATA2[2];
  assign n102 = DATA1[4];
  assign n111 = DATA1[17];
  assign n123 = DATA1[3];
  assign n125 = DATA1[1];
  assign n126 = DATA1[0];
  assign n127 = DATA2[1];
  assign n128 = DATA1[2];
  assign n129 = DATA1[5];
  assign n130 = DATA1[8];
  assign n131 = DATA1[10];
  assign n132 = DATA1[11];
  assign n133 = DATA1[12];
  assign n134 = DATA1[13];
  assign n135 = DATA1[15];
  assign n136 = DATA1[16];
  assign n137 = DATA1[20];
  assign n138 = DATA1[21];
  assign n139 = DATA1[22];
  assign n140 = DATA1[23];
  assign n141 = DATA1[24];
  assign n142 = DATA1[25];
  assign n143 = DATA1[26];
  assign n144 = DATA1[28];

  RCA_GEN_NBIT32 adder4 ( .A({DATA1[31], n91, DATA1[29], n171, n89, n170, n169, 
        n168, n167, n166, n165, n164, DATA1[19:18], n111, n163, n162, 
        DATA1[14], n161, n160, n159, n158, n74, n130, n157, n156, n155, n102, 
        n154, n128, n125, n126}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0}), .Ci(1'b0), .S(return_address) );
  SHIFTER_GENERIC_N32 shifter ( .A({DATA1[31], n91, DATA1[29], n171, n89, n170, 
        n169, n168, n167, n166, n165, n164, DATA1[19:18], n111, n163, n162, 
        DATA1[14], n161, n160, n159, n158, n74, n130, n157, n156, n155, n102, 
        n154, n149, n150, n153}), .B({DATA2[4:3], n152, n151, n58}), 
        .LOGIC_ARITH(ShiftOpCode[2]), .LEFT_RIGHT(ShiftOpCode[1]), 
        .SHIFT_ROTATE(ShiftOpCode[0]), .OUTPUT(shift_out) );
  operatore_logic_REG_SIZE32 logic_operations ( .A({DATA1[31], n91, DATA1[29], 
        n171, n89, n170, n169, n168, n167, n166, n165, n164, DATA1[19:18], 
        n111, n163, n162, DATA1[14], n161, n160, n159, n158, n74, n130, n157, 
        n156, n155, n102, n154, n149, n150, n153}), .B({DATA2[31:3], n152, 
        n151, n58}), .OUT_LOGIC_AND(AND_OUT), .OUT_LOGIC_OR(OR_OUT), 
        .OUT_LOGIC_XOR(XOR_OUT) );
  p4_adder_N32_N_carry4 adder_sub ( .A({DATA1[31], n91, DATA1[29], n171, n89, 
        n170, n169, n168, n167, n166, n165, n164, DATA1[19:18], n111, n163, 
        n162, DATA1[14], n161, n160, n159, n158, n74, n130, n157, n156, n155, 
        n102, n154, n149, n150, n153}), .B({DATA2[31:3], n152, n151, n58}), 
        .Cin(Add_subn), .SUM(add_sub_out) );
  compare_N32 comp ( .num1({DATA1[31], n91, DATA1[29], n171, n89, n170, n169, 
        n168, n167, n166, n165, n164, DATA1[19:18], n111, n163, n162, 
        DATA1[14], n161, n160, n159, n158, n74, n130, n157, n156, n155, n102, 
        n154, n128, n148, n153}), .num2({DATA2[31:3], n152, n127, n58}), 
        .equal(comp_eq), .greater(comp_greater) );
  MUX_2to1_n32 mux_comp ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1}), .S(sel_mux_comp_out), 
        .Y(comp_out) );
  MUX_6to1_n32 mux_alu_out ( .A(add_sub_out), .B(AND_OUT), .C(OR_OUT), .D(
        XOR_OUT), .E(comp_out), .F(shift_out), .S(AluOpCode), .Y(OUTALU) );
  BUF_X1 U3 ( .A(n127), .Z(n151) );
  INV_X1 U4 ( .A(CompareOpCode[2]), .ZN(n146) );
  INV_X1 U5 ( .A(CompareOpCode[3]), .ZN(n147) );
  CLKBUF_X2 U6 ( .A(n138), .Z(n165) );
  CLKBUF_X2 U7 ( .A(n140), .Z(n167) );
  OAI22_X1 U8 ( .A1(n146), .A2(comp_eq), .B1(n5), .B2(n147), .ZN(CompBranch)
         );
  BUF_X4 U9 ( .A(n129), .Z(n155) );
  INV_X1 U10 ( .A(comp_eq), .ZN(n5) );
  NAND2_X1 U11 ( .A1(n3), .A2(n4), .ZN(sel_mux_comp_out) );
  OAI21_X1 U12 ( .B1(comp_eq), .B2(comp_greater), .A(CompareOpCode[1]), .ZN(n4) );
  NAND2_X1 U13 ( .A1(CompareOpCode[0]), .A2(n5), .ZN(n3) );
  BUF_X2 U14 ( .A(n139), .Z(n166) );
  BUF_X2 U15 ( .A(n137), .Z(n164) );
  BUF_X2 U16 ( .A(n134), .Z(n161) );
  BUF_X2 U17 ( .A(n143), .Z(n170) );
  BUF_X2 U18 ( .A(n135), .Z(n162) );
  BUF_X2 U19 ( .A(n133), .Z(n160) );
  BUF_X2 U20 ( .A(n132), .Z(n159) );
  BUF_X2 U21 ( .A(n131), .Z(n158) );
  BUF_X2 U22 ( .A(n71), .Z(n156) );
  BUF_X2 U23 ( .A(n136), .Z(n163) );
  BUF_X2 U24 ( .A(n141), .Z(n168) );
  BUF_X2 U25 ( .A(n142), .Z(n169) );
  BUF_X2 U26 ( .A(n144), .Z(n171) );
  BUF_X2 U27 ( .A(n72), .Z(n157) );
  CLKBUF_X1 U28 ( .A(n125), .Z(n148) );
  BUF_X4 U29 ( .A(n123), .Z(n154) );
  CLKBUF_X1 U30 ( .A(n128), .Z(n149) );
  CLKBUF_X1 U31 ( .A(n148), .Z(n150) );
  CLKBUF_X1 U32 ( .A(n126), .Z(n153) );
  CLKBUF_X3 U33 ( .A(n100), .Z(n152) );
endmodule


module mux21_N32_3 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n118, n119, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136;

  INV_X2 U63 ( .A(n66), .ZN(Y[0]) );
  BUF_X1 U1 ( .A(n124), .Z(n132) );
  INV_X1 U2 ( .A(n41), .ZN(Y[3]) );
  BUF_X1 U3 ( .A(n125), .Z(n136) );
  NOR2_X1 U4 ( .A1(n121), .A2(n123), .ZN(n118) );
  NOR2_X1 U5 ( .A1(n122), .A2(n127), .ZN(n119) );
  OR2_X1 U6 ( .A1(n118), .A2(n119), .ZN(Y[1]) );
  INV_X1 U7 ( .A(A[1]), .ZN(n121) );
  INV_X1 U8 ( .A(B[1]), .ZN(n122) );
  INV_X1 U9 ( .A(n136), .ZN(n127) );
  CLKBUF_X1 U10 ( .A(n125), .Z(n135) );
  CLKBUF_X1 U11 ( .A(n125), .Z(n134) );
  INV_X1 U12 ( .A(n136), .ZN(n126) );
  BUF_X1 U13 ( .A(n123), .Z(n129) );
  CLKBUF_X1 U14 ( .A(n123), .Z(n128) );
  CLKBUF_X1 U15 ( .A(n124), .Z(n133) );
  CLKBUF_X1 U16 ( .A(n124), .Z(n131) );
  CLKBUF_X1 U17 ( .A(n123), .Z(n130) );
  AOI22_X1 U18 ( .A1(A[3]), .A2(n127), .B1(B[3]), .B2(n129), .ZN(n41) );
  INV_X1 U19 ( .A(n39), .ZN(Y[5]) );
  AOI22_X1 U20 ( .A1(A[5]), .A2(n127), .B1(B[5]), .B2(n128), .ZN(n39) );
  INV_X1 U21 ( .A(n38), .ZN(Y[6]) );
  AOI22_X1 U22 ( .A1(A[6]), .A2(n127), .B1(B[6]), .B2(n128), .ZN(n38) );
  INV_X1 U23 ( .A(n44), .ZN(Y[2]) );
  AOI22_X1 U24 ( .A1(A[2]), .A2(n126), .B1(B[2]), .B2(n129), .ZN(n44) );
  INV_X1 U25 ( .A(n64), .ZN(Y[11]) );
  AOI22_X1 U26 ( .A1(A[11]), .A2(n126), .B1(B[11]), .B2(n135), .ZN(n64) );
  AOI22_X1 U27 ( .A1(A[0]), .A2(n127), .B1(B[0]), .B2(n135), .ZN(n66) );
  INV_X1 U28 ( .A(n63), .ZN(Y[12]) );
  AOI22_X1 U29 ( .A1(A[12]), .A2(n126), .B1(B[12]), .B2(n134), .ZN(n63) );
  INV_X1 U30 ( .A(n62), .ZN(Y[13]) );
  AOI22_X1 U31 ( .A1(A[13]), .A2(n126), .B1(B[13]), .B2(n134), .ZN(n62) );
  INV_X1 U32 ( .A(n61), .ZN(Y[14]) );
  AOI22_X1 U33 ( .A1(A[14]), .A2(n126), .B1(B[14]), .B2(n134), .ZN(n61) );
  INV_X1 U34 ( .A(n60), .ZN(Y[15]) );
  AOI22_X1 U35 ( .A1(A[15]), .A2(n126), .B1(B[15]), .B2(n134), .ZN(n60) );
  INV_X1 U36 ( .A(n59), .ZN(Y[16]) );
  AOI22_X1 U37 ( .A1(A[16]), .A2(n126), .B1(B[16]), .B2(n133), .ZN(n59) );
  INV_X1 U38 ( .A(n57), .ZN(Y[18]) );
  AOI22_X1 U39 ( .A1(A[18]), .A2(n127), .B1(B[18]), .B2(n133), .ZN(n57) );
  INV_X1 U40 ( .A(n51), .ZN(Y[23]) );
  AOI22_X1 U41 ( .A1(A[23]), .A2(n126), .B1(B[23]), .B2(n131), .ZN(n51) );
  INV_X1 U42 ( .A(n49), .ZN(Y[25]) );
  AOI22_X1 U43 ( .A1(A[25]), .A2(n126), .B1(B[25]), .B2(n131), .ZN(n49) );
  INV_X1 U44 ( .A(n47), .ZN(Y[27]) );
  AOI22_X1 U45 ( .A1(A[27]), .A2(n126), .B1(B[27]), .B2(n130), .ZN(n47) );
  INV_X1 U46 ( .A(n50), .ZN(Y[24]) );
  AOI22_X1 U47 ( .A1(A[24]), .A2(n126), .B1(B[24]), .B2(n131), .ZN(n50) );
  INV_X1 U48 ( .A(n46), .ZN(Y[28]) );
  AOI22_X1 U49 ( .A1(A[28]), .A2(n126), .B1(B[28]), .B2(n130), .ZN(n46) );
  INV_X1 U50 ( .A(n58), .ZN(Y[17]) );
  AOI22_X1 U51 ( .A1(A[17]), .A2(n126), .B1(B[17]), .B2(n133), .ZN(n58) );
  INV_X1 U52 ( .A(n43), .ZN(Y[30]) );
  AOI22_X1 U53 ( .A1(A[30]), .A2(n126), .B1(B[30]), .B2(n132), .ZN(n43) );
  INV_X1 U54 ( .A(n54), .ZN(Y[20]) );
  AOI22_X1 U55 ( .A1(A[20]), .A2(n126), .B1(B[20]), .B2(n132), .ZN(n54) );
  INV_X1 U56 ( .A(n48), .ZN(Y[26]) );
  AOI22_X1 U57 ( .A1(A[26]), .A2(n126), .B1(B[26]), .B2(n130), .ZN(n48) );
  INV_X1 U58 ( .A(n56), .ZN(Y[19]) );
  AOI22_X1 U59 ( .A1(A[19]), .A2(n126), .B1(B[19]), .B2(n133), .ZN(n56) );
  INV_X1 U60 ( .A(n45), .ZN(Y[29]) );
  AOI22_X1 U61 ( .A1(A[29]), .A2(n126), .B1(B[29]), .B2(n130), .ZN(n45) );
  INV_X1 U62 ( .A(n53), .ZN(Y[21]) );
  AOI22_X1 U64 ( .A1(A[21]), .A2(n126), .B1(B[21]), .B2(n132), .ZN(n53) );
  INV_X1 U65 ( .A(n65), .ZN(Y[10]) );
  AOI22_X1 U66 ( .A1(A[10]), .A2(n126), .B1(B[10]), .B2(n135), .ZN(n65) );
  INV_X1 U67 ( .A(n52), .ZN(Y[22]) );
  AOI22_X1 U68 ( .A1(A[22]), .A2(n126), .B1(B[22]), .B2(n131), .ZN(n52) );
  INV_X1 U69 ( .A(n34), .ZN(Y[9]) );
  AOI22_X1 U70 ( .A1(A[9]), .A2(n127), .B1(n135), .B2(B[9]), .ZN(n34) );
  INV_X1 U71 ( .A(n37), .ZN(Y[7]) );
  AOI22_X1 U72 ( .A1(A[7]), .A2(n127), .B1(B[7]), .B2(n128), .ZN(n37) );
  INV_X1 U73 ( .A(n36), .ZN(Y[8]) );
  AOI22_X1 U74 ( .A1(A[8]), .A2(n127), .B1(B[8]), .B2(n128), .ZN(n36) );
  INV_X1 U75 ( .A(n40), .ZN(Y[4]) );
  AOI22_X1 U76 ( .A1(A[4]), .A2(n127), .B1(B[4]), .B2(n129), .ZN(n40) );
  INV_X1 U77 ( .A(n42), .ZN(Y[31]) );
  AOI22_X1 U78 ( .A1(A[31]), .A2(n127), .B1(B[31]), .B2(n129), .ZN(n42) );
  CLKBUF_X1 U79 ( .A(SEL), .Z(n123) );
  CLKBUF_X1 U80 ( .A(SEL), .Z(n124) );
  BUF_X1 U81 ( .A(SEL), .Z(n125) );
endmodule


module mux21_N32_4 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   net77012, net167276, n36, n37, n38, n39, n40, n43, n44, n45, n46, n47,
         n48, n49, n50, n51, n52, n53, n54, n55, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n99, n100, n101, n103, n105, n106, n107, n109,
         n110, n111, n112, n113, n114, n115, n116, n117;
  assign net77012 = SEL;
  assign Y[0] = net167276;

  INV_X1 U1 ( .A(A[4]), .ZN(n105) );
  INV_X1 U2 ( .A(B[4]), .ZN(n106) );
  INV_X1 U3 ( .A(n58), .ZN(Y[18]) );
  BUF_X1 U4 ( .A(net77012), .Z(n110) );
  CLKBUF_X1 U5 ( .A(net77012), .Z(n99) );
  CLKBUF_X1 U6 ( .A(n113), .Z(n117) );
  BUF_X2 U7 ( .A(n99), .Z(n113) );
  NOR2_X1 U8 ( .A1(n107), .A2(n112), .ZN(n100) );
  OR2_X1 U9 ( .A1(n100), .A2(n101), .ZN(Y[3]) );
  AND2_X1 U10 ( .A1(A[3]), .A2(n112), .ZN(n101) );
  BUF_X1 U11 ( .A(n99), .Z(n103) );
  OAI22_X4 U12 ( .A1(n105), .A2(n113), .B1(n106), .B2(n112), .ZN(Y[4]) );
  INV_X1 U13 ( .A(n110), .ZN(n111) );
  INV_X1 U14 ( .A(B[3]), .ZN(n107) );
  MUX2_X1 U15 ( .A(A[0]), .B(B[0]), .S(net77012), .Z(net167276) );
  MUX2_X1 U16 ( .A(A[1]), .B(B[1]), .S(n110), .Z(Y[1]) );
  INV_X1 U17 ( .A(n53), .ZN(Y[22]) );
  INV_X1 U18 ( .A(n55), .ZN(Y[20]) );
  INV_X1 U19 ( .A(n57), .ZN(Y[19]) );
  INV_X1 U20 ( .A(n63), .ZN(Y[13]) );
  INV_X1 U21 ( .A(n49), .ZN(Y[26]) );
  INV_X1 U22 ( .A(n61), .ZN(Y[15]) );
  INV_X1 U23 ( .A(n62), .ZN(Y[14]) );
  INV_X1 U24 ( .A(n37), .ZN(Y[8]) );
  INV_X1 U25 ( .A(n43), .ZN(Y[31]) );
  INV_X1 U26 ( .A(n64), .ZN(Y[12]) );
  INV_X1 U27 ( .A(n54), .ZN(Y[21]) );
  INV_X1 U28 ( .A(n52), .ZN(Y[23]) );
  INV_X1 U29 ( .A(n65), .ZN(Y[11]) );
  INV_X1 U30 ( .A(n59), .ZN(Y[17]) );
  INV_X1 U31 ( .A(n48), .ZN(Y[27]) );
  INV_X1 U32 ( .A(n44), .ZN(Y[30]) );
  INV_X1 U33 ( .A(n36), .ZN(Y[9]) );
  INV_X1 U34 ( .A(n66), .ZN(Y[10]) );
  INV_X1 U35 ( .A(n39), .ZN(Y[6]) );
  INV_X1 U36 ( .A(n60), .ZN(Y[16]) );
  INV_X1 U37 ( .A(n46), .ZN(Y[29]) );
  INV_X1 U38 ( .A(n40), .ZN(Y[5]) );
  INV_X1 U39 ( .A(n51), .ZN(Y[24]) );
  INV_X1 U40 ( .A(n50), .ZN(Y[25]) );
  INV_X1 U41 ( .A(n47), .ZN(Y[28]) );
  INV_X1 U42 ( .A(n38), .ZN(Y[7]) );
  BUF_X1 U43 ( .A(n103), .Z(n114) );
  INV_X1 U44 ( .A(net77012), .ZN(n112) );
  INV_X1 U45 ( .A(n113), .ZN(n109) );
  CLKBUF_X1 U46 ( .A(n99), .Z(n116) );
  INV_X1 U47 ( .A(n45), .ZN(Y[2]) );
  CLKBUF_X1 U48 ( .A(n99), .Z(n115) );
  AOI22_X1 U49 ( .A1(A[31]), .A2(n109), .B1(B[31]), .B2(n113), .ZN(n43) );
  AOI22_X1 U50 ( .A1(A[30]), .A2(n109), .B1(B[30]), .B2(n114), .ZN(n44) );
  AOI22_X1 U51 ( .A1(A[27]), .A2(n109), .B1(B[27]), .B2(n116), .ZN(n48) );
  AOI22_X1 U52 ( .A1(A[26]), .A2(n109), .B1(B[26]), .B2(n114), .ZN(n49) );
  AOI22_X1 U53 ( .A1(A[23]), .A2(n109), .B1(B[23]), .B2(n114), .ZN(n52) );
  AOI22_X1 U54 ( .A1(A[22]), .A2(n109), .B1(B[22]), .B2(n113), .ZN(n53) );
  AOI22_X1 U55 ( .A1(A[20]), .A2(n109), .B1(B[20]), .B2(n116), .ZN(n55) );
  AOI22_X1 U56 ( .A1(A[17]), .A2(n109), .B1(B[17]), .B2(n103), .ZN(n59) );
  AOI22_X1 U57 ( .A1(A[15]), .A2(n109), .B1(B[15]), .B2(n117), .ZN(n61) );
  AOI22_X1 U58 ( .A1(A[13]), .A2(n109), .B1(B[13]), .B2(n117), .ZN(n63) );
  AOI22_X1 U59 ( .A1(A[11]), .A2(n109), .B1(B[11]), .B2(n115), .ZN(n65) );
  AOI22_X1 U60 ( .A1(A[29]), .A2(n111), .B1(B[29]), .B2(n103), .ZN(n46) );
  AOI22_X1 U61 ( .A1(A[28]), .A2(n111), .B1(B[28]), .B2(n115), .ZN(n47) );
  AOI22_X1 U62 ( .A1(A[25]), .A2(n111), .B1(B[25]), .B2(n114), .ZN(n50) );
  AOI22_X1 U63 ( .A1(A[24]), .A2(n111), .B1(B[24]), .B2(n114), .ZN(n51) );
  AOI22_X1 U64 ( .A1(A[21]), .A2(n111), .B1(B[21]), .B2(n115), .ZN(n54) );
  AOI22_X1 U65 ( .A1(A[19]), .A2(n111), .B1(B[19]), .B2(n103), .ZN(n57) );
  AOI22_X1 U66 ( .A1(A[18]), .A2(n111), .B1(B[18]), .B2(n113), .ZN(n58) );
  AOI22_X1 U67 ( .A1(A[16]), .A2(n111), .B1(B[16]), .B2(n117), .ZN(n60) );
  AOI22_X1 U68 ( .A1(A[14]), .A2(n111), .B1(B[14]), .B2(n117), .ZN(n62) );
  AOI22_X1 U69 ( .A1(A[12]), .A2(n111), .B1(B[12]), .B2(n116), .ZN(n64) );
  AOI22_X1 U70 ( .A1(A[10]), .A2(n111), .B1(B[10]), .B2(n103), .ZN(n66) );
  AOI22_X1 U71 ( .A1(A[2]), .A2(n112), .B1(B[2]), .B2(n110), .ZN(n45) );
  AOI22_X1 U72 ( .A1(A[9]), .A2(n111), .B1(B[9]), .B2(n115), .ZN(n36) );
  AOI22_X1 U73 ( .A1(A[8]), .A2(n111), .B1(B[8]), .B2(n116), .ZN(n37) );
  AOI22_X1 U74 ( .A1(A[7]), .A2(n111), .B1(B[7]), .B2(n115), .ZN(n38) );
  AOI22_X1 U75 ( .A1(A[6]), .A2(n111), .B1(B[6]), .B2(n116), .ZN(n39) );
  AOI22_X1 U76 ( .A1(A[5]), .A2(n111), .B1(B[5]), .B2(n103), .ZN(n40) );
endmodule


module registro_N5_0 ( data, enable, clock, clear, Q );
  input [4:0] data;
  output [4:0] Q;
  input enable, clock, clear;
  wire   n11, n12, n13, n14, n15, net44619, net44620, net44621, net44622,
         net44623, n1, n2, n3, n4, n5;
  tri   enable;

  DFFR_X1 \Q_reg[4]  ( .D(n15), .CK(clock), .RN(clear), .Q(Q[4]), .QN(net44623) );
  DFFR_X1 \Q_reg[3]  ( .D(n14), .CK(clock), .RN(clear), .Q(Q[3]), .QN(net44622) );
  DFFR_X1 \Q_reg[2]  ( .D(n13), .CK(clock), .RN(clear), .Q(Q[2]), .QN(net44621) );
  DFFR_X1 \Q_reg[1]  ( .D(n12), .CK(clock), .RN(clear), .Q(Q[1]), .QN(net44620) );
  DFFR_X1 \Q_reg[0]  ( .D(n11), .CK(clock), .RN(clear), .Q(Q[0]), .QN(net44619) );
  OAI21_X1 U2 ( .B1(net44619), .B2(enable), .A(n5), .ZN(n11) );
  NAND2_X1 U3 ( .A1(data[0]), .A2(enable), .ZN(n5) );
  OAI21_X1 U4 ( .B1(net44620), .B2(enable), .A(n4), .ZN(n12) );
  NAND2_X1 U5 ( .A1(data[1]), .A2(enable), .ZN(n4) );
  OAI21_X1 U6 ( .B1(net44621), .B2(enable), .A(n3), .ZN(n13) );
  NAND2_X1 U7 ( .A1(data[2]), .A2(enable), .ZN(n3) );
  OAI21_X1 U8 ( .B1(net44622), .B2(enable), .A(n2), .ZN(n14) );
  NAND2_X1 U9 ( .A1(data[3]), .A2(enable), .ZN(n2) );
  OAI21_X1 U10 ( .B1(net44623), .B2(enable), .A(n1), .ZN(n15) );
  NAND2_X1 U11 ( .A1(enable), .A2(data[4]), .ZN(n1) );
endmodule


module registro_N17 ( data, enable, clock, clear, Q );
  input [16:0] data;
  output [16:0] Q;
  input enable, clock, clear;
  wire   n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, net44602, net44603, net44604, net44605, net44606,
         net44607, net44608, net44609, net44610, net44611, net44612, net44613,
         net44614, net44615, net44616, net44617, net44618, n59, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n60, n61,
         n62, n63, n64;
  assign n59 = clear;

  DFFR_X1 \Q_reg[16]  ( .D(n51), .CK(clock), .RN(n60), .Q(Q[16]), .QN(net44618) );
  DFFR_X1 \Q_reg[15]  ( .D(n50), .CK(clock), .RN(n60), .Q(Q[15]), .QN(net44617) );
  DFFR_X1 \Q_reg[14]  ( .D(n49), .CK(clock), .RN(n60), .Q(Q[14]), .QN(net44616) );
  DFFR_X1 \Q_reg[13]  ( .D(n48), .CK(clock), .RN(n60), .Q(Q[13]), .QN(net44615) );
  DFFR_X1 \Q_reg[12]  ( .D(n47), .CK(clock), .RN(n60), .Q(Q[12]), .QN(net44614) );
  DFFR_X1 \Q_reg[11]  ( .D(n46), .CK(clock), .RN(n61), .Q(Q[11]), .QN(net44613) );
  DFFR_X1 \Q_reg[10]  ( .D(n45), .CK(clock), .RN(n61), .Q(Q[10]), .QN(net44612) );
  DFFR_X1 \Q_reg[9]  ( .D(n44), .CK(clock), .RN(n61), .Q(Q[9]), .QN(net44611)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n43), .CK(clock), .RN(n61), .Q(Q[8]), .QN(net44610)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n42), .CK(clock), .RN(n60), .Q(Q[7]), .QN(net44609)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n41), .CK(clock), .RN(n60), .Q(Q[6]), .QN(net44608)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n40), .CK(clock), .RN(n60), .Q(Q[5]), .QN(net44607)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n39), .CK(clock), .RN(n61), .Q(Q[4]), .QN(net44606)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n38), .CK(clock), .RN(n60), .Q(Q[3]), .QN(net44605)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n37), .CK(clock), .RN(n60), .Q(Q[2]), .QN(net44604)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n36), .CK(clock), .RN(n61), .Q(Q[1]), .QN(net44603)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n35), .CK(clock), .RN(n60), .Q(Q[0]), .QN(net44602)
         );
  BUF_X1 U2 ( .A(enable), .Z(n62) );
  BUF_X1 U3 ( .A(enable), .Z(n63) );
  BUF_X1 U4 ( .A(enable), .Z(n64) );
  BUF_X1 U5 ( .A(n59), .Z(n60) );
  BUF_X1 U6 ( .A(n59), .Z(n61) );
  OAI21_X1 U7 ( .B1(net44605), .B2(n63), .A(n14), .ZN(n38) );
  NAND2_X1 U8 ( .A1(data[3]), .A2(n63), .ZN(n14) );
  OAI21_X1 U9 ( .B1(net44606), .B2(n63), .A(n13), .ZN(n39) );
  NAND2_X1 U10 ( .A1(data[4]), .A2(n63), .ZN(n13) );
  OAI21_X1 U11 ( .B1(net44607), .B2(n63), .A(n12), .ZN(n40) );
  NAND2_X1 U12 ( .A1(data[5]), .A2(n62), .ZN(n12) );
  OAI21_X1 U13 ( .B1(net44608), .B2(n63), .A(n11), .ZN(n41) );
  NAND2_X1 U14 ( .A1(data[6]), .A2(n62), .ZN(n11) );
  OAI21_X1 U15 ( .B1(net44609), .B2(n63), .A(n10), .ZN(n42) );
  NAND2_X1 U16 ( .A1(data[7]), .A2(n62), .ZN(n10) );
  OAI21_X1 U17 ( .B1(net44610), .B2(n63), .A(n9), .ZN(n43) );
  NAND2_X1 U18 ( .A1(data[8]), .A2(n62), .ZN(n9) );
  OAI21_X1 U19 ( .B1(net44611), .B2(n63), .A(n8), .ZN(n44) );
  NAND2_X1 U20 ( .A1(data[9]), .A2(n62), .ZN(n8) );
  OAI21_X1 U21 ( .B1(net44612), .B2(n63), .A(n7), .ZN(n45) );
  NAND2_X1 U22 ( .A1(data[10]), .A2(n62), .ZN(n7) );
  OAI21_X1 U23 ( .B1(net44602), .B2(n64), .A(n17), .ZN(n35) );
  NAND2_X1 U24 ( .A1(data[0]), .A2(n62), .ZN(n17) );
  OAI21_X1 U25 ( .B1(net44603), .B2(n64), .A(n16), .ZN(n36) );
  NAND2_X1 U26 ( .A1(data[1]), .A2(n63), .ZN(n16) );
  OAI21_X1 U27 ( .B1(net44604), .B2(n64), .A(n15), .ZN(n37) );
  NAND2_X1 U28 ( .A1(data[2]), .A2(n63), .ZN(n15) );
  OAI21_X1 U29 ( .B1(net44613), .B2(n64), .A(n6), .ZN(n46) );
  NAND2_X1 U30 ( .A1(data[11]), .A2(n62), .ZN(n6) );
  OAI21_X1 U31 ( .B1(net44614), .B2(n64), .A(n5), .ZN(n47) );
  NAND2_X1 U32 ( .A1(data[12]), .A2(n62), .ZN(n5) );
  OAI21_X1 U33 ( .B1(net44615), .B2(n64), .A(n4), .ZN(n48) );
  NAND2_X1 U34 ( .A1(data[13]), .A2(n62), .ZN(n4) );
  OAI21_X1 U35 ( .B1(net44616), .B2(n64), .A(n3), .ZN(n49) );
  NAND2_X1 U36 ( .A1(data[14]), .A2(n62), .ZN(n3) );
  OAI21_X1 U37 ( .B1(net44617), .B2(n64), .A(n2), .ZN(n50) );
  NAND2_X1 U38 ( .A1(data[15]), .A2(n62), .ZN(n2) );
  OAI21_X1 U39 ( .B1(net44618), .B2(n64), .A(n1), .ZN(n51) );
  NAND2_X1 U40 ( .A1(n64), .A2(data[16]), .ZN(n1) );
endmodule


module registro_N32_6 ( data, enable, clock, clear, Q );
  input [31:0] data;
  output [31:0] Q;
  input enable, clock, clear;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net44624, net44625, net44626, net44627, net44628, net44629,
         net44630, net44631, net44632, net44633, net44634, net44635, net44636,
         net44637, net44638, net44639, net44640, net44641, net44642, net44643,
         net44644, net44645, net44646, net44647, net44648, net44649, net44650,
         net44651, net44652, net44653, net44654, net44655, n111, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n112, n113, n114;
  tri   enable;
  assign n111 = clear;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(clock), .RN(n114), .Q(Q[31]), .QN(net44655) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(clock), .RN(n114), .Q(Q[30]), .QN(net44654) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(clock), .RN(n114), .Q(Q[29]), .QN(net44653) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(clock), .RN(n114), .Q(Q[28]), .QN(net44652) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(clock), .RN(n114), .Q(Q[27]), .QN(net44651) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(clock), .RN(n114), .Q(Q[26]), .QN(net44650) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(clock), .RN(n114), .Q(Q[25]), .QN(net44649) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(clock), .RN(n114), .Q(Q[24]), .QN(net44648) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(clock), .RN(n114), .Q(Q[23]), .QN(net44647) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(clock), .RN(n114), .Q(Q[22]), .QN(
        net44646) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(clock), .RN(n112), .Q(Q[21]), .QN(
        net44645) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(clock), .RN(n112), .Q(Q[20]), .QN(
        net44644) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(clock), .RN(n112), .Q(Q[19]), .QN(
        net44643) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(clock), .RN(n112), .Q(Q[18]), .QN(
        net44642) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(clock), .RN(n112), .Q(Q[17]), .QN(
        net44641) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(clock), .RN(n112), .Q(Q[16]), .QN(
        net44640) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(clock), .RN(n112), .Q(Q[15]), .QN(
        net44639) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(clock), .RN(n112), .Q(Q[14]), .QN(
        net44638) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(clock), .RN(n112), .Q(Q[13]), .QN(
        net44637) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(clock), .RN(n112), .Q(Q[12]), .QN(
        net44636) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(clock), .RN(n112), .Q(Q[11]), .QN(
        net44635) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(clock), .RN(n113), .Q(Q[10]), .QN(
        net44634) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(clock), .RN(n113), .Q(Q[9]), .QN(net44633)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(clock), .RN(n113), .Q(Q[8]), .QN(net44632)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(clock), .RN(n113), .Q(Q[7]), .QN(net44631)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(clock), .RN(n113), .Q(Q[6]), .QN(net44630)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(clock), .RN(n113), .Q(Q[5]), .QN(net44629)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(clock), .RN(n113), .Q(Q[4]), .QN(net44628)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(clock), .RN(n113), .Q(Q[3]), .QN(net44627)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(clock), .RN(n113), .Q(Q[2]), .QN(net44626)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(clock), .RN(n113), .Q(Q[1]), .QN(net44625)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(clock), .RN(n113), .Q(Q[0]), .QN(net44624)
         );
  BUF_X1 U2 ( .A(n111), .Z(n113) );
  BUF_X1 U3 ( .A(n111), .Z(n112) );
  BUF_X1 U4 ( .A(n111), .Z(n114) );
  OAI21_X1 U5 ( .B1(net44647), .B2(enable), .A(n33), .ZN(n9) );
  NAND2_X1 U6 ( .A1(enable), .A2(data[23]), .ZN(n33) );
  OAI21_X1 U7 ( .B1(net44624), .B2(enable), .A(n39), .ZN(n32) );
  NAND2_X1 U8 ( .A1(data[0]), .A2(enable), .ZN(n39) );
  OAI21_X1 U9 ( .B1(net44625), .B2(enable), .A(n40), .ZN(n31) );
  NAND2_X1 U10 ( .A1(data[1]), .A2(enable), .ZN(n40) );
  OAI21_X1 U11 ( .B1(net44626), .B2(enable), .A(n41), .ZN(n30) );
  NAND2_X1 U12 ( .A1(data[2]), .A2(enable), .ZN(n41) );
  OAI21_X1 U13 ( .B1(net44627), .B2(enable), .A(n43), .ZN(n29) );
  NAND2_X1 U14 ( .A1(data[3]), .A2(enable), .ZN(n43) );
  OAI21_X1 U15 ( .B1(net44628), .B2(enable), .A(n44), .ZN(n28) );
  NAND2_X1 U16 ( .A1(data[4]), .A2(enable), .ZN(n44) );
  OAI21_X1 U17 ( .B1(net44629), .B2(enable), .A(n45), .ZN(n27) );
  NAND2_X1 U18 ( .A1(data[5]), .A2(enable), .ZN(n45) );
  OAI21_X1 U19 ( .B1(net44630), .B2(enable), .A(n46), .ZN(n26) );
  NAND2_X1 U20 ( .A1(data[6]), .A2(enable), .ZN(n46) );
  OAI21_X1 U21 ( .B1(net44631), .B2(enable), .A(n47), .ZN(n25) );
  NAND2_X1 U22 ( .A1(data[7]), .A2(enable), .ZN(n47) );
  OAI21_X1 U23 ( .B1(net44632), .B2(enable), .A(n48), .ZN(n24) );
  NAND2_X1 U24 ( .A1(data[8]), .A2(enable), .ZN(n48) );
  OAI21_X1 U25 ( .B1(net44633), .B2(enable), .A(n49), .ZN(n23) );
  NAND2_X1 U26 ( .A1(data[9]), .A2(enable), .ZN(n49) );
  OAI21_X1 U27 ( .B1(net44634), .B2(enable), .A(n50), .ZN(n22) );
  NAND2_X1 U28 ( .A1(data[10]), .A2(enable), .ZN(n50) );
  OAI21_X1 U29 ( .B1(net44635), .B2(enable), .A(n51), .ZN(n21) );
  NAND2_X1 U30 ( .A1(data[11]), .A2(enable), .ZN(n51) );
  OAI21_X1 U31 ( .B1(net44636), .B2(enable), .A(n52), .ZN(n20) );
  NAND2_X1 U32 ( .A1(data[12]), .A2(enable), .ZN(n52) );
  OAI21_X1 U33 ( .B1(net44637), .B2(enable), .A(n54), .ZN(n19) );
  NAND2_X1 U34 ( .A1(data[13]), .A2(enable), .ZN(n54) );
  OAI21_X1 U35 ( .B1(net44638), .B2(enable), .A(n55), .ZN(n18) );
  NAND2_X1 U36 ( .A1(data[14]), .A2(enable), .ZN(n55) );
  OAI21_X1 U37 ( .B1(net44639), .B2(enable), .A(n56), .ZN(n17) );
  NAND2_X1 U38 ( .A1(data[15]), .A2(enable), .ZN(n56) );
  OAI21_X1 U39 ( .B1(net44640), .B2(enable), .A(n57), .ZN(n16) );
  NAND2_X1 U40 ( .A1(data[16]), .A2(enable), .ZN(n57) );
  OAI21_X1 U41 ( .B1(net44641), .B2(enable), .A(n58), .ZN(n15) );
  NAND2_X1 U42 ( .A1(data[17]), .A2(enable), .ZN(n58) );
  OAI21_X1 U43 ( .B1(net44642), .B2(enable), .A(n59), .ZN(n14) );
  NAND2_X1 U44 ( .A1(data[18]), .A2(enable), .ZN(n59) );
  OAI21_X1 U45 ( .B1(net44643), .B2(enable), .A(n60), .ZN(n13) );
  NAND2_X1 U46 ( .A1(data[19]), .A2(enable), .ZN(n60) );
  OAI21_X1 U47 ( .B1(net44644), .B2(enable), .A(n61), .ZN(n12) );
  NAND2_X1 U48 ( .A1(data[20]), .A2(enable), .ZN(n61) );
  OAI21_X1 U49 ( .B1(net44645), .B2(enable), .A(n62), .ZN(n11) );
  NAND2_X1 U50 ( .A1(data[21]), .A2(enable), .ZN(n62) );
  OAI21_X1 U51 ( .B1(net44646), .B2(enable), .A(n63), .ZN(n10) );
  NAND2_X1 U52 ( .A1(data[22]), .A2(enable), .ZN(n63) );
  OAI21_X1 U53 ( .B1(net44648), .B2(enable), .A(n34), .ZN(n8) );
  NAND2_X1 U54 ( .A1(data[24]), .A2(enable), .ZN(n34) );
  OAI21_X1 U55 ( .B1(net44649), .B2(enable), .A(n35), .ZN(n7) );
  NAND2_X1 U56 ( .A1(data[25]), .A2(enable), .ZN(n35) );
  OAI21_X1 U57 ( .B1(net44650), .B2(enable), .A(n36), .ZN(n6) );
  NAND2_X1 U58 ( .A1(data[26]), .A2(enable), .ZN(n36) );
  OAI21_X1 U59 ( .B1(net44651), .B2(enable), .A(n37), .ZN(n5) );
  NAND2_X1 U60 ( .A1(data[27]), .A2(enable), .ZN(n37) );
  OAI21_X1 U61 ( .B1(net44652), .B2(enable), .A(n38), .ZN(n4) );
  NAND2_X1 U62 ( .A1(data[28]), .A2(enable), .ZN(n38) );
  OAI21_X1 U63 ( .B1(net44653), .B2(enable), .A(n42), .ZN(n3) );
  NAND2_X1 U64 ( .A1(data[29]), .A2(enable), .ZN(n42) );
  OAI21_X1 U65 ( .B1(net44654), .B2(enable), .A(n53), .ZN(n2) );
  NAND2_X1 U66 ( .A1(data[30]), .A2(enable), .ZN(n53) );
  OAI21_X1 U67 ( .B1(net44655), .B2(enable), .A(n64), .ZN(n1) );
  NAND2_X1 U68 ( .A1(data[31]), .A2(enable), .ZN(n64) );
endmodule


module registro_N32_7 ( data, enable, clock, clear, Q );
  input [31:0] data;
  output [31:0] Q;
  input enable, clock, clear;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net44624, net44625, net44626, net44627, net44628, net44629,
         net44630, net44631, net44632, net44633, net44634, net44635, net44636,
         net44637, net44638, net44639, net44640, net44641, net44642, net44643,
         net44644, net44645, net44646, net44647, net44648, net44649, net44650,
         net44651, net44652, net44653, net44654, net44655, n141, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n142, n143, n144, n145, n146, n147, n148, n149, n150;
  assign n141 = clear;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(clock), .RN(n144), .Q(Q[31]), .QN(net44655) );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(clock), .RN(n144), .Q(Q[30]), .QN(net44654) );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(clock), .RN(n144), .Q(Q[29]), .QN(net44653) );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(clock), .RN(n144), .Q(Q[28]), .QN(net44652) );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(clock), .RN(n144), .Q(Q[27]), .QN(net44651) );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(clock), .RN(n144), .Q(Q[26]), .QN(net44650) );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(clock), .RN(n144), .Q(Q[25]), .QN(net44649) );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(clock), .RN(n144), .Q(Q[24]), .QN(net44648) );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(clock), .RN(n144), .Q(Q[23]), .QN(net44647) );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(clock), .RN(n144), .Q(Q[22]), .QN(
        net44646) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(clock), .RN(n142), .Q(Q[21]), .QN(
        net44645) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(clock), .RN(n142), .Q(Q[20]), .QN(
        net44644) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(clock), .RN(n142), .Q(Q[19]), .QN(
        net44643) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(clock), .RN(n142), .Q(Q[18]), .QN(
        net44642) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(clock), .RN(n142), .Q(Q[17]), .QN(
        net44641) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(clock), .RN(n142), .Q(Q[16]), .QN(
        net44640) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(clock), .RN(n142), .Q(Q[15]), .QN(
        net44639) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(clock), .RN(n142), .Q(Q[14]), .QN(
        net44638) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(clock), .RN(n142), .Q(Q[13]), .QN(
        net44637) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(clock), .RN(n142), .Q(Q[12]), .QN(
        net44636) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(clock), .RN(n142), .Q(Q[11]), .QN(
        net44635) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(clock), .RN(n143), .Q(Q[10]), .QN(
        net44634) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(clock), .RN(n143), .Q(Q[9]), .QN(net44633)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(clock), .RN(n143), .Q(Q[8]), .QN(net44632)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(clock), .RN(n143), .Q(Q[7]), .QN(net44631)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(clock), .RN(n143), .Q(Q[6]), .QN(net44630)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(clock), .RN(n143), .Q(Q[5]), .QN(net44629)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(clock), .RN(n143), .Q(Q[4]), .QN(net44628)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(clock), .RN(n143), .Q(Q[3]), .QN(net44627)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(clock), .RN(n143), .Q(Q[2]), .QN(net44626)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(clock), .RN(n143), .Q(Q[1]), .QN(net44625)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(clock), .RN(n143), .Q(Q[0]), .QN(net44624)
         );
  BUF_X1 U2 ( .A(n141), .Z(n143) );
  BUF_X1 U3 ( .A(n141), .Z(n142) );
  BUF_X1 U4 ( .A(n141), .Z(n144) );
  OAI21_X1 U5 ( .B1(net44624), .B2(n148), .A(n39), .ZN(n32) );
  NAND2_X1 U6 ( .A1(data[0]), .A2(n146), .ZN(n39) );
  OAI21_X1 U7 ( .B1(net44625), .B2(n147), .A(n40), .ZN(n31) );
  NAND2_X1 U8 ( .A1(data[1]), .A2(n146), .ZN(n40) );
  OAI21_X1 U9 ( .B1(net44626), .B2(n148), .A(n41), .ZN(n30) );
  NAND2_X1 U10 ( .A1(data[2]), .A2(n146), .ZN(n41) );
  OAI21_X1 U11 ( .B1(net44627), .B2(n148), .A(n43), .ZN(n29) );
  NAND2_X1 U12 ( .A1(data[3]), .A2(n146), .ZN(n43) );
  OAI21_X1 U13 ( .B1(net44634), .B2(n149), .A(n50), .ZN(n22) );
  NAND2_X1 U14 ( .A1(data[10]), .A2(n146), .ZN(n50) );
  OAI21_X1 U15 ( .B1(net44635), .B2(n149), .A(n51), .ZN(n21) );
  NAND2_X1 U16 ( .A1(data[11]), .A2(n146), .ZN(n51) );
  OAI21_X1 U17 ( .B1(net44636), .B2(n149), .A(n52), .ZN(n20) );
  NAND2_X1 U18 ( .A1(data[12]), .A2(n146), .ZN(n52) );
  OAI21_X1 U19 ( .B1(net44637), .B2(n149), .A(n54), .ZN(n19) );
  NAND2_X1 U20 ( .A1(data[13]), .A2(n146), .ZN(n54) );
  OAI21_X1 U21 ( .B1(net44638), .B2(n149), .A(n55), .ZN(n18) );
  NAND2_X1 U22 ( .A1(data[14]), .A2(n146), .ZN(n55) );
  OAI21_X1 U23 ( .B1(net44639), .B2(n149), .A(n56), .ZN(n17) );
  NAND2_X1 U24 ( .A1(data[15]), .A2(n146), .ZN(n56) );
  OAI21_X1 U25 ( .B1(net44640), .B2(n149), .A(n57), .ZN(n16) );
  NAND2_X1 U26 ( .A1(data[16]), .A2(n145), .ZN(n57) );
  OAI21_X1 U27 ( .B1(net44641), .B2(n149), .A(n58), .ZN(n15) );
  NAND2_X1 U28 ( .A1(data[17]), .A2(n145), .ZN(n58) );
  OAI21_X1 U29 ( .B1(net44642), .B2(n149), .A(n59), .ZN(n14) );
  NAND2_X1 U30 ( .A1(data[18]), .A2(n145), .ZN(n59) );
  OAI21_X1 U31 ( .B1(net44643), .B2(n149), .A(n60), .ZN(n13) );
  NAND2_X1 U32 ( .A1(data[19]), .A2(n145), .ZN(n60) );
  OAI21_X1 U33 ( .B1(net44644), .B2(n150), .A(n61), .ZN(n12) );
  NAND2_X1 U34 ( .A1(data[20]), .A2(n145), .ZN(n61) );
  OAI21_X1 U35 ( .B1(net44645), .B2(n150), .A(n62), .ZN(n11) );
  NAND2_X1 U36 ( .A1(data[21]), .A2(n145), .ZN(n62) );
  OAI21_X1 U37 ( .B1(net44646), .B2(n150), .A(n63), .ZN(n10) );
  NAND2_X1 U38 ( .A1(data[22]), .A2(n145), .ZN(n63) );
  OAI21_X1 U39 ( .B1(net44648), .B2(n147), .A(n34), .ZN(n8) );
  NAND2_X1 U40 ( .A1(data[24]), .A2(n145), .ZN(n34) );
  OAI21_X1 U41 ( .B1(net44649), .B2(n147), .A(n35), .ZN(n7) );
  NAND2_X1 U42 ( .A1(data[25]), .A2(n145), .ZN(n35) );
  OAI21_X1 U43 ( .B1(net44650), .B2(n148), .A(n36), .ZN(n6) );
  NAND2_X1 U44 ( .A1(data[26]), .A2(n145), .ZN(n36) );
  OAI21_X1 U45 ( .B1(net44651), .B2(n147), .A(n37), .ZN(n5) );
  NAND2_X1 U46 ( .A1(data[27]), .A2(n145), .ZN(n37) );
  OAI21_X1 U47 ( .B1(net44652), .B2(n147), .A(n38), .ZN(n4) );
  NAND2_X1 U48 ( .A1(data[28]), .A2(n146), .ZN(n38) );
  OAI21_X1 U49 ( .B1(net44654), .B2(n149), .A(n53), .ZN(n2) );
  NAND2_X1 U50 ( .A1(data[30]), .A2(n146), .ZN(n53) );
  OAI21_X1 U51 ( .B1(net44655), .B2(n148), .A(n64), .ZN(n1) );
  NAND2_X1 U52 ( .A1(data[31]), .A2(n145), .ZN(n64) );
  OAI21_X1 U53 ( .B1(net44628), .B2(n148), .A(n44), .ZN(n28) );
  NAND2_X1 U54 ( .A1(data[4]), .A2(n147), .ZN(n44) );
  OAI21_X1 U55 ( .B1(net44629), .B2(n148), .A(n45), .ZN(n27) );
  NAND2_X1 U56 ( .A1(data[5]), .A2(n147), .ZN(n45) );
  OAI21_X1 U57 ( .B1(net44630), .B2(n148), .A(n46), .ZN(n26) );
  NAND2_X1 U58 ( .A1(data[6]), .A2(n147), .ZN(n46) );
  OAI21_X1 U59 ( .B1(net44631), .B2(n148), .A(n47), .ZN(n25) );
  NAND2_X1 U60 ( .A1(data[7]), .A2(n147), .ZN(n47) );
  OAI21_X1 U61 ( .B1(net44632), .B2(n148), .A(n48), .ZN(n24) );
  NAND2_X1 U62 ( .A1(data[8]), .A2(n147), .ZN(n48) );
  OAI21_X1 U63 ( .B1(net44633), .B2(n149), .A(n49), .ZN(n23) );
  NAND2_X1 U64 ( .A1(data[9]), .A2(n147), .ZN(n49) );
  OAI21_X1 U65 ( .B1(net44653), .B2(n148), .A(n42), .ZN(n3) );
  NAND2_X1 U66 ( .A1(data[29]), .A2(n147), .ZN(n42) );
  OAI21_X1 U67 ( .B1(net44647), .B2(n148), .A(n33), .ZN(n9) );
  NAND2_X1 U68 ( .A1(n150), .A2(data[23]), .ZN(n33) );
  CLKBUF_X1 U69 ( .A(enable), .Z(n145) );
  CLKBUF_X1 U70 ( .A(enable), .Z(n146) );
  CLKBUF_X1 U71 ( .A(enable), .Z(n147) );
  CLKBUF_X1 U72 ( .A(enable), .Z(n148) );
  CLKBUF_X1 U73 ( .A(enable), .Z(n149) );
  CLKBUF_X1 U74 ( .A(enable), .Z(n150) );
endmodule


module registro_N32_8 ( data, enable, clock, clear, Q );
  input [31:0] data;
  output [31:0] Q;
  input enable, clock, clear;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, net44624, net44625, net44626, net44627, net44628, net44629,
         net44630, net44631, net44632, net44633, net44634, net44635, net44636,
         net44637, net44638, net44639, net44640, net44641, net44642, net44643,
         net44644, net44645, net44646, net44647, net44648, net44649, net44650,
         net44651, net44652, net44653, net44654, net44655, n79, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n80, n81, n82;
  tri   enable;
  assign n79 = clear;

  DFFR_X1 \Q_reg[31]  ( .D(n1), .CK(clock), .RN(n82), .Q(Q[31]), .QN(net44655)
         );
  DFFR_X1 \Q_reg[30]  ( .D(n2), .CK(clock), .RN(n82), .Q(Q[30]), .QN(net44654)
         );
  DFFR_X1 \Q_reg[29]  ( .D(n3), .CK(clock), .RN(n82), .Q(Q[29]), .QN(net44653)
         );
  DFFR_X1 \Q_reg[28]  ( .D(n4), .CK(clock), .RN(n82), .Q(Q[28]), .QN(net44652)
         );
  DFFR_X1 \Q_reg[27]  ( .D(n5), .CK(clock), .RN(n82), .Q(Q[27]), .QN(net44651)
         );
  DFFR_X1 \Q_reg[26]  ( .D(n6), .CK(clock), .RN(n82), .Q(Q[26]), .QN(net44650)
         );
  DFFR_X1 \Q_reg[25]  ( .D(n7), .CK(clock), .RN(n82), .Q(Q[25]), .QN(net44649)
         );
  DFFR_X1 \Q_reg[24]  ( .D(n8), .CK(clock), .RN(n82), .Q(Q[24]), .QN(net44648)
         );
  DFFR_X1 \Q_reg[23]  ( .D(n9), .CK(clock), .RN(n82), .Q(Q[23]), .QN(net44647)
         );
  DFFR_X1 \Q_reg[22]  ( .D(n10), .CK(clock), .RN(n82), .Q(Q[22]), .QN(net44646) );
  DFFR_X1 \Q_reg[21]  ( .D(n11), .CK(clock), .RN(n80), .Q(Q[21]), .QN(net44645) );
  DFFR_X1 \Q_reg[20]  ( .D(n12), .CK(clock), .RN(n80), .Q(Q[20]), .QN(net44644) );
  DFFR_X1 \Q_reg[19]  ( .D(n13), .CK(clock), .RN(n80), .Q(Q[19]), .QN(net44643) );
  DFFR_X1 \Q_reg[18]  ( .D(n14), .CK(clock), .RN(n80), .Q(Q[18]), .QN(net44642) );
  DFFR_X1 \Q_reg[17]  ( .D(n15), .CK(clock), .RN(n80), .Q(Q[17]), .QN(net44641) );
  DFFR_X1 \Q_reg[16]  ( .D(n16), .CK(clock), .RN(n80), .Q(Q[16]), .QN(net44640) );
  DFFR_X1 \Q_reg[15]  ( .D(n17), .CK(clock), .RN(n80), .Q(Q[15]), .QN(net44639) );
  DFFR_X1 \Q_reg[14]  ( .D(n18), .CK(clock), .RN(n80), .Q(Q[14]), .QN(net44638) );
  DFFR_X1 \Q_reg[13]  ( .D(n19), .CK(clock), .RN(n80), .Q(Q[13]), .QN(net44637) );
  DFFR_X1 \Q_reg[12]  ( .D(n20), .CK(clock), .RN(n80), .Q(Q[12]), .QN(net44636) );
  DFFR_X1 \Q_reg[11]  ( .D(n21), .CK(clock), .RN(n80), .Q(Q[11]), .QN(net44635) );
  DFFR_X1 \Q_reg[10]  ( .D(n22), .CK(clock), .RN(n81), .Q(Q[10]), .QN(net44634) );
  DFFR_X1 \Q_reg[9]  ( .D(n23), .CK(clock), .RN(n81), .Q(Q[9]), .QN(net44633)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n24), .CK(clock), .RN(n81), .Q(Q[8]), .QN(net44632)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n25), .CK(clock), .RN(n81), .Q(Q[7]), .QN(net44631)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n26), .CK(clock), .RN(n81), .Q(Q[6]), .QN(net44630)
         );
  DFFR_X1 \Q_reg[5]  ( .D(n27), .CK(clock), .RN(n81), .Q(Q[5]), .QN(net44629)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n28), .CK(clock), .RN(n81), .Q(Q[4]), .QN(net44628)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n29), .CK(clock), .RN(n81), .Q(Q[3]), .QN(net44627)
         );
  DFFR_X1 \Q_reg[2]  ( .D(n30), .CK(clock), .RN(n81), .Q(Q[2]), .QN(net44626)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n31), .CK(clock), .RN(n81), .Q(Q[1]), .QN(net44625)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n32), .CK(clock), .RN(n81), .Q(Q[0]), .QN(net44624)
         );
  BUF_X1 U2 ( .A(n79), .Z(n81) );
  BUF_X1 U3 ( .A(n79), .Z(n80) );
  BUF_X1 U4 ( .A(n79), .Z(n82) );
  OAI21_X1 U5 ( .B1(net44647), .B2(enable), .A(n33), .ZN(n9) );
  NAND2_X1 U6 ( .A1(enable), .A2(data[23]), .ZN(n33) );
  OAI21_X1 U7 ( .B1(net44624), .B2(enable), .A(n39), .ZN(n32) );
  NAND2_X1 U8 ( .A1(data[0]), .A2(enable), .ZN(n39) );
  OAI21_X1 U9 ( .B1(net44625), .B2(enable), .A(n40), .ZN(n31) );
  NAND2_X1 U10 ( .A1(data[1]), .A2(enable), .ZN(n40) );
  OAI21_X1 U11 ( .B1(net44626), .B2(enable), .A(n41), .ZN(n30) );
  NAND2_X1 U12 ( .A1(data[2]), .A2(enable), .ZN(n41) );
  OAI21_X1 U13 ( .B1(net44627), .B2(enable), .A(n43), .ZN(n29) );
  NAND2_X1 U14 ( .A1(data[3]), .A2(enable), .ZN(n43) );
  OAI21_X1 U15 ( .B1(net44628), .B2(enable), .A(n44), .ZN(n28) );
  NAND2_X1 U16 ( .A1(data[4]), .A2(enable), .ZN(n44) );
  OAI21_X1 U17 ( .B1(net44629), .B2(enable), .A(n45), .ZN(n27) );
  NAND2_X1 U18 ( .A1(data[5]), .A2(enable), .ZN(n45) );
  OAI21_X1 U19 ( .B1(net44630), .B2(enable), .A(n46), .ZN(n26) );
  NAND2_X1 U20 ( .A1(data[6]), .A2(enable), .ZN(n46) );
  OAI21_X1 U21 ( .B1(net44631), .B2(enable), .A(n47), .ZN(n25) );
  NAND2_X1 U22 ( .A1(data[7]), .A2(enable), .ZN(n47) );
  OAI21_X1 U23 ( .B1(net44632), .B2(enable), .A(n48), .ZN(n24) );
  NAND2_X1 U24 ( .A1(data[8]), .A2(enable), .ZN(n48) );
  OAI21_X1 U25 ( .B1(net44633), .B2(enable), .A(n49), .ZN(n23) );
  NAND2_X1 U26 ( .A1(data[9]), .A2(enable), .ZN(n49) );
  OAI21_X1 U27 ( .B1(net44634), .B2(enable), .A(n50), .ZN(n22) );
  NAND2_X1 U28 ( .A1(data[10]), .A2(enable), .ZN(n50) );
  OAI21_X1 U29 ( .B1(net44635), .B2(enable), .A(n51), .ZN(n21) );
  NAND2_X1 U30 ( .A1(data[11]), .A2(enable), .ZN(n51) );
  OAI21_X1 U31 ( .B1(net44636), .B2(enable), .A(n52), .ZN(n20) );
  NAND2_X1 U32 ( .A1(data[12]), .A2(enable), .ZN(n52) );
  OAI21_X1 U33 ( .B1(net44637), .B2(enable), .A(n54), .ZN(n19) );
  NAND2_X1 U34 ( .A1(data[13]), .A2(enable), .ZN(n54) );
  OAI21_X1 U35 ( .B1(net44638), .B2(enable), .A(n55), .ZN(n18) );
  NAND2_X1 U36 ( .A1(data[14]), .A2(enable), .ZN(n55) );
  OAI21_X1 U37 ( .B1(net44639), .B2(enable), .A(n56), .ZN(n17) );
  NAND2_X1 U38 ( .A1(data[15]), .A2(enable), .ZN(n56) );
  OAI21_X1 U39 ( .B1(net44640), .B2(enable), .A(n57), .ZN(n16) );
  NAND2_X1 U40 ( .A1(data[16]), .A2(enable), .ZN(n57) );
  OAI21_X1 U41 ( .B1(net44641), .B2(enable), .A(n58), .ZN(n15) );
  NAND2_X1 U42 ( .A1(data[17]), .A2(enable), .ZN(n58) );
  OAI21_X1 U43 ( .B1(net44642), .B2(enable), .A(n59), .ZN(n14) );
  NAND2_X1 U44 ( .A1(data[18]), .A2(enable), .ZN(n59) );
  OAI21_X1 U45 ( .B1(net44643), .B2(enable), .A(n60), .ZN(n13) );
  NAND2_X1 U46 ( .A1(data[19]), .A2(enable), .ZN(n60) );
  OAI21_X1 U47 ( .B1(net44644), .B2(enable), .A(n61), .ZN(n12) );
  NAND2_X1 U48 ( .A1(data[20]), .A2(enable), .ZN(n61) );
  OAI21_X1 U49 ( .B1(net44645), .B2(enable), .A(n62), .ZN(n11) );
  NAND2_X1 U50 ( .A1(data[21]), .A2(enable), .ZN(n62) );
  OAI21_X1 U51 ( .B1(net44646), .B2(enable), .A(n63), .ZN(n10) );
  NAND2_X1 U52 ( .A1(data[22]), .A2(enable), .ZN(n63) );
  OAI21_X1 U53 ( .B1(net44648), .B2(enable), .A(n34), .ZN(n8) );
  NAND2_X1 U54 ( .A1(data[24]), .A2(enable), .ZN(n34) );
  OAI21_X1 U55 ( .B1(net44649), .B2(enable), .A(n35), .ZN(n7) );
  NAND2_X1 U56 ( .A1(data[25]), .A2(enable), .ZN(n35) );
  OAI21_X1 U57 ( .B1(net44650), .B2(enable), .A(n36), .ZN(n6) );
  NAND2_X1 U58 ( .A1(data[26]), .A2(enable), .ZN(n36) );
  OAI21_X1 U59 ( .B1(net44651), .B2(enable), .A(n37), .ZN(n5) );
  NAND2_X1 U60 ( .A1(data[27]), .A2(enable), .ZN(n37) );
  OAI21_X1 U61 ( .B1(net44652), .B2(enable), .A(n38), .ZN(n4) );
  NAND2_X1 U62 ( .A1(data[28]), .A2(enable), .ZN(n38) );
  OAI21_X1 U63 ( .B1(net44653), .B2(enable), .A(n42), .ZN(n3) );
  NAND2_X1 U64 ( .A1(data[29]), .A2(enable), .ZN(n42) );
  OAI21_X1 U65 ( .B1(net44654), .B2(enable), .A(n53), .ZN(n2) );
  NAND2_X1 U66 ( .A1(data[30]), .A2(enable), .ZN(n53) );
  OAI21_X1 U67 ( .B1(net44655), .B2(enable), .A(n64), .ZN(n1) );
  NAND2_X1 U68 ( .A1(data[31]), .A2(enable), .ZN(n64) );
endmodule


module registro_N32_0 ( data, enable, clock, clear, Q );
  input [31:0] data;
  output [31:0] Q;
  input enable, clock, clear;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, net44570, net44571, net44572, net44573, net44574,
         net44575, net44576, net44577, net44578, net44579, net44580, net44581,
         net44582, net44583, net44584, net44585, net44586, net44587, net44588,
         net44589, net44590, net44591, net44592, net44593, net44594, net44595,
         net44596, net44597, net44598, net44599, net44600, net44601, n47, n1,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n48, n49, n50;
  tri   enable;
  assign n47 = clear;

  DFFR_X1 \Q_reg[31]  ( .D(n96), .CK(clock), .RN(n50), .Q(Q[31]), .QN(net44601) );
  DFFR_X1 \Q_reg[29]  ( .D(n94), .CK(clock), .RN(n50), .Q(Q[29]), .QN(net44599) );
  DFFR_X1 \Q_reg[28]  ( .D(n93), .CK(clock), .RN(n50), .Q(Q[28]), .QN(net44598) );
  DFFR_X1 \Q_reg[26]  ( .D(n91), .CK(clock), .RN(n48), .Q(Q[26]), .QN(net44596) );
  DFFR_X1 \Q_reg[25]  ( .D(n90), .CK(clock), .RN(n49), .Q(Q[25]), .QN(net44595) );
  DFFR_X1 \Q_reg[24]  ( .D(n89), .CK(clock), .RN(n49), .Q(Q[24]), .QN(net44594) );
  DFFR_X1 \Q_reg[22]  ( .D(n87), .CK(clock), .RN(n48), .Q(Q[22]), .QN(net44592) );
  DFFR_X1 \Q_reg[20]  ( .D(n85), .CK(clock), .RN(n50), .Q(Q[20]), .QN(net44590) );
  DFFR_X1 \Q_reg[19]  ( .D(n84), .CK(clock), .RN(n48), .Q(Q[19]), .QN(net44589) );
  DFFR_X1 \Q_reg[18]  ( .D(n83), .CK(clock), .RN(n50), .Q(Q[18]), .QN(net44588) );
  DFFR_X1 \Q_reg[16]  ( .D(n81), .CK(clock), .RN(n49), .Q(Q[16]), .QN(net44586) );
  DFFR_X1 \Q_reg[15]  ( .D(n80), .CK(clock), .RN(n49), .Q(Q[15]), .QN(net44585) );
  DFFR_X1 \Q_reg[14]  ( .D(n79), .CK(clock), .RN(n49), .Q(Q[14]), .QN(net44584) );
  DFFR_X1 \Q_reg[10]  ( .D(n75), .CK(clock), .RN(n50), .Q(Q[10]), .QN(net44580) );
  DFFR_X1 \Q_reg[2]  ( .D(n67), .CK(clock), .RN(n48), .Q(Q[2]), .QN(net44572)
         );
  DFFR_X1 \Q_reg[1]  ( .D(n66), .CK(clock), .RN(n48), .Q(Q[1]), .QN(net44571)
         );
  DFFR_X1 \Q_reg[0]  ( .D(n65), .CK(clock), .RN(n48), .Q(Q[0]), .QN(net44570)
         );
  DFFR_X1 \Q_reg[13]  ( .D(n78), .CK(clock), .RN(n48), .Q(Q[13]), .QN(net44583) );
  DFFR_X1 \Q_reg[12]  ( .D(n77), .CK(clock), .RN(n48), .Q(Q[12]), .QN(net44582) );
  DFFR_X1 \Q_reg[11]  ( .D(n76), .CK(clock), .RN(n50), .Q(Q[11]), .QN(net44581) );
  DFFR_X1 \Q_reg[9]  ( .D(n74), .CK(clock), .RN(n49), .Q(Q[9]), .QN(net44579)
         );
  DFFR_X1 \Q_reg[7]  ( .D(n72), .CK(clock), .RN(n49), .Q(Q[7]), .QN(net44577)
         );
  DFFR_X1 \Q_reg[6]  ( .D(n71), .CK(clock), .RN(n49), .Q(Q[6]), .QN(net44576)
         );
  DFFR_X1 \Q_reg[4]  ( .D(n69), .CK(clock), .RN(n49), .Q(Q[4]), .QN(net44574)
         );
  DFFR_X1 \Q_reg[8]  ( .D(n73), .CK(clock), .RN(n49), .Q(Q[8]), .QN(net44578)
         );
  DFFR_X1 \Q_reg[3]  ( .D(n68), .CK(clock), .RN(n48), .Q(Q[3]), .QN(net44573)
         );
  DFFR_X1 \Q_reg[17]  ( .D(n82), .CK(clock), .RN(n50), .Q(Q[17]), .QN(net44587) );
  DFFR_X1 \Q_reg[23]  ( .D(n88), .CK(clock), .RN(n49), .Q(Q[23]), .QN(net44593) );
  DFFR_X1 \Q_reg[27]  ( .D(n92), .CK(clock), .RN(n50), .Q(Q[27]), .QN(net44597) );
  DFFR_X1 \Q_reg[30]  ( .D(n95), .CK(clock), .RN(n50), .Q(Q[30]), .QN(net44600) );
  DFFR_X1 \Q_reg[21]  ( .D(n86), .CK(clock), .RN(n48), .Q(Q[21]), .QN(net44591) );
  DFFR_X1 \Q_reg[5]  ( .D(n70), .CK(clock), .RN(n48), .Q(Q[5]), .QN(net44575)
         );
  BUF_X1 U2 ( .A(n47), .Z(n49) );
  BUF_X1 U3 ( .A(n47), .Z(n48) );
  BUF_X1 U4 ( .A(n47), .Z(n50) );
  OAI21_X1 U5 ( .B1(net44601), .B2(enable), .A(n1), .ZN(n96) );
  NAND2_X1 U6 ( .A1(enable), .A2(data[31]), .ZN(n1) );
  OAI21_X1 U7 ( .B1(net44591), .B2(enable), .A(n11), .ZN(n86) );
  NAND2_X1 U8 ( .A1(data[21]), .A2(enable), .ZN(n11) );
  OAI21_X1 U9 ( .B1(net44600), .B2(enable), .A(n2), .ZN(n95) );
  NAND2_X1 U10 ( .A1(data[30]), .A2(enable), .ZN(n2) );
  OAI21_X1 U11 ( .B1(net44597), .B2(enable), .A(n5), .ZN(n92) );
  NAND2_X1 U12 ( .A1(data[27]), .A2(enable), .ZN(n5) );
  OAI21_X1 U13 ( .B1(net44575), .B2(enable), .A(n27), .ZN(n70) );
  NAND2_X1 U14 ( .A1(data[5]), .A2(enable), .ZN(n27) );
  OAI21_X1 U15 ( .B1(net44573), .B2(enable), .A(n29), .ZN(n68) );
  NAND2_X1 U16 ( .A1(data[3]), .A2(enable), .ZN(n29) );
  OAI21_X1 U17 ( .B1(net44578), .B2(enable), .A(n24), .ZN(n73) );
  NAND2_X1 U18 ( .A1(data[8]), .A2(enable), .ZN(n24) );
  OAI21_X1 U19 ( .B1(net44593), .B2(enable), .A(n9), .ZN(n88) );
  NAND2_X1 U20 ( .A1(data[23]), .A2(enable), .ZN(n9) );
  OAI21_X1 U21 ( .B1(net44574), .B2(enable), .A(n28), .ZN(n69) );
  NAND2_X1 U22 ( .A1(data[4]), .A2(enable), .ZN(n28) );
  OAI21_X1 U23 ( .B1(net44576), .B2(enable), .A(n26), .ZN(n71) );
  NAND2_X1 U24 ( .A1(data[6]), .A2(enable), .ZN(n26) );
  OAI21_X1 U25 ( .B1(net44577), .B2(enable), .A(n25), .ZN(n72) );
  NAND2_X1 U26 ( .A1(data[7]), .A2(enable), .ZN(n25) );
  OAI21_X1 U27 ( .B1(net44579), .B2(enable), .A(n23), .ZN(n74) );
  NAND2_X1 U28 ( .A1(data[9]), .A2(enable), .ZN(n23) );
  OAI21_X1 U29 ( .B1(net44581), .B2(enable), .A(n21), .ZN(n76) );
  NAND2_X1 U30 ( .A1(data[11]), .A2(enable), .ZN(n21) );
  OAI21_X1 U31 ( .B1(net44582), .B2(enable), .A(n20), .ZN(n77) );
  NAND2_X1 U32 ( .A1(data[12]), .A2(enable), .ZN(n20) );
  OAI21_X1 U33 ( .B1(net44583), .B2(enable), .A(n19), .ZN(n78) );
  NAND2_X1 U34 ( .A1(data[13]), .A2(enable), .ZN(n19) );
  OAI21_X1 U35 ( .B1(net44570), .B2(enable), .A(n32), .ZN(n65) );
  NAND2_X1 U36 ( .A1(data[0]), .A2(enable), .ZN(n32) );
  OAI21_X1 U37 ( .B1(net44571), .B2(enable), .A(n31), .ZN(n66) );
  NAND2_X1 U38 ( .A1(data[1]), .A2(enable), .ZN(n31) );
  OAI21_X1 U39 ( .B1(net44572), .B2(enable), .A(n30), .ZN(n67) );
  NAND2_X1 U40 ( .A1(data[2]), .A2(enable), .ZN(n30) );
  OAI21_X1 U41 ( .B1(net44580), .B2(enable), .A(n22), .ZN(n75) );
  NAND2_X1 U42 ( .A1(data[10]), .A2(enable), .ZN(n22) );
  OAI21_X1 U43 ( .B1(net44584), .B2(enable), .A(n18), .ZN(n79) );
  NAND2_X1 U44 ( .A1(data[14]), .A2(enable), .ZN(n18) );
  OAI21_X1 U45 ( .B1(net44585), .B2(enable), .A(n17), .ZN(n80) );
  NAND2_X1 U46 ( .A1(data[15]), .A2(enable), .ZN(n17) );
  OAI21_X1 U47 ( .B1(net44586), .B2(enable), .A(n16), .ZN(n81) );
  NAND2_X1 U48 ( .A1(data[16]), .A2(enable), .ZN(n16) );
  OAI21_X1 U49 ( .B1(net44587), .B2(enable), .A(n15), .ZN(n82) );
  NAND2_X1 U50 ( .A1(data[17]), .A2(enable), .ZN(n15) );
  OAI21_X1 U51 ( .B1(net44588), .B2(enable), .A(n14), .ZN(n83) );
  NAND2_X1 U52 ( .A1(data[18]), .A2(enable), .ZN(n14) );
  OAI21_X1 U53 ( .B1(net44589), .B2(enable), .A(n13), .ZN(n84) );
  NAND2_X1 U54 ( .A1(data[19]), .A2(enable), .ZN(n13) );
  OAI21_X1 U55 ( .B1(net44590), .B2(enable), .A(n12), .ZN(n85) );
  NAND2_X1 U56 ( .A1(data[20]), .A2(enable), .ZN(n12) );
  OAI21_X1 U57 ( .B1(net44592), .B2(enable), .A(n10), .ZN(n87) );
  NAND2_X1 U58 ( .A1(data[22]), .A2(enable), .ZN(n10) );
  OAI21_X1 U59 ( .B1(net44594), .B2(enable), .A(n8), .ZN(n89) );
  NAND2_X1 U60 ( .A1(data[24]), .A2(enable), .ZN(n8) );
  OAI21_X1 U61 ( .B1(net44595), .B2(enable), .A(n7), .ZN(n90) );
  NAND2_X1 U62 ( .A1(data[25]), .A2(enable), .ZN(n7) );
  OAI21_X1 U63 ( .B1(net44596), .B2(enable), .A(n6), .ZN(n91) );
  NAND2_X1 U64 ( .A1(data[26]), .A2(enable), .ZN(n6) );
  OAI21_X1 U65 ( .B1(net44598), .B2(enable), .A(n4), .ZN(n93) );
  NAND2_X1 U66 ( .A1(data[28]), .A2(enable), .ZN(n4) );
  OAI21_X1 U67 ( .B1(net44599), .B2(enable), .A(n3), .ZN(n94) );
  NAND2_X1 U68 ( .A1(data[29]), .A2(enable), .ZN(n3) );
endmodule


module SIG_EXT_BITS32 ( EXT_UNSIGNED, EXT_FOR_J, S_IN, S_OUT );
  input [31:0] S_IN;
  output [31:0] S_OUT;
  input EXT_UNSIGNED, EXT_FOR_J;
  wire   \S_OUT[26] , \S_IN[15] , \S_IN[14] , \S_IN[13] , \S_IN[12] ,
         \S_IN[11] , \S_IN[10] , \S_IN[9] , \S_IN[8] , \S_IN[7] , \S_IN[6] ,
         \S_IN[5] , \S_IN[4] , \S_IN[3] , \S_IN[2] , \S_IN[1] , \S_IN[0] , n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17;
  assign S_OUT[31] = \S_OUT[26] ;
  assign S_OUT[30] = \S_OUT[26] ;
  assign S_OUT[29] = \S_OUT[26] ;
  assign S_OUT[28] = \S_OUT[26] ;
  assign S_OUT[27] = \S_OUT[26] ;
  assign S_OUT[26] = \S_OUT[26] ;
  assign S_OUT[15] = \S_IN[15] ;
  assign \S_IN[15]  = S_IN[15];
  assign S_OUT[14] = \S_IN[14] ;
  assign \S_IN[14]  = S_IN[14];
  assign S_OUT[13] = \S_IN[13] ;
  assign \S_IN[13]  = S_IN[13];
  assign S_OUT[12] = \S_IN[12] ;
  assign \S_IN[12]  = S_IN[12];
  assign S_OUT[11] = \S_IN[11] ;
  assign \S_IN[11]  = S_IN[11];
  assign S_OUT[10] = \S_IN[10] ;
  assign \S_IN[10]  = S_IN[10];
  assign S_OUT[9] = \S_IN[9] ;
  assign \S_IN[9]  = S_IN[9];
  assign S_OUT[8] = \S_IN[8] ;
  assign \S_IN[8]  = S_IN[8];
  assign S_OUT[7] = \S_IN[7] ;
  assign \S_IN[7]  = S_IN[7];
  assign S_OUT[6] = \S_IN[6] ;
  assign \S_IN[6]  = S_IN[6];
  assign S_OUT[5] = \S_IN[5] ;
  assign \S_IN[5]  = S_IN[5];
  assign S_OUT[4] = \S_IN[4] ;
  assign \S_IN[4]  = S_IN[4];
  assign S_OUT[3] = \S_IN[3] ;
  assign \S_IN[3]  = S_IN[3];
  assign S_OUT[2] = \S_IN[2] ;
  assign \S_IN[2]  = S_IN[2];
  assign S_OUT[1] = \S_IN[1] ;
  assign \S_IN[1]  = S_IN[1];
  assign S_OUT[0] = \S_IN[0] ;
  assign \S_IN[0]  = S_IN[0];

  NAND3_X1 U25 ( .A1(EXT_FOR_J), .A2(n6), .A3(S_IN[25]), .ZN(n5) );
  NAND2_X1 U2 ( .A1(n4), .A2(n10), .ZN(S_OUT[23]) );
  NAND2_X1 U3 ( .A1(S_IN[23]), .A2(EXT_FOR_J), .ZN(n10) );
  NAND2_X1 U4 ( .A1(n4), .A2(n17), .ZN(S_OUT[16]) );
  NAND2_X1 U5 ( .A1(S_IN[16]), .A2(EXT_FOR_J), .ZN(n17) );
  NAND2_X1 U6 ( .A1(n4), .A2(n16), .ZN(S_OUT[17]) );
  NAND2_X1 U7 ( .A1(S_IN[17]), .A2(EXT_FOR_J), .ZN(n16) );
  NAND2_X1 U8 ( .A1(n4), .A2(n15), .ZN(S_OUT[18]) );
  NAND2_X1 U9 ( .A1(S_IN[18]), .A2(EXT_FOR_J), .ZN(n15) );
  NAND2_X1 U10 ( .A1(n4), .A2(n14), .ZN(S_OUT[19]) );
  NAND2_X1 U11 ( .A1(S_IN[19]), .A2(EXT_FOR_J), .ZN(n14) );
  NAND2_X1 U12 ( .A1(n4), .A2(n13), .ZN(S_OUT[20]) );
  NAND2_X1 U13 ( .A1(S_IN[20]), .A2(EXT_FOR_J), .ZN(n13) );
  NAND2_X1 U14 ( .A1(n4), .A2(n12), .ZN(S_OUT[21]) );
  NAND2_X1 U15 ( .A1(S_IN[21]), .A2(EXT_FOR_J), .ZN(n12) );
  NAND2_X1 U16 ( .A1(n4), .A2(n11), .ZN(S_OUT[22]) );
  NAND2_X1 U17 ( .A1(S_IN[22]), .A2(EXT_FOR_J), .ZN(n11) );
  NAND2_X1 U18 ( .A1(n4), .A2(n9), .ZN(S_OUT[24]) );
  NAND2_X1 U19 ( .A1(S_IN[24]), .A2(EXT_FOR_J), .ZN(n9) );
  OAI21_X1 U20 ( .B1(n7), .B2(n8), .A(n4), .ZN(S_OUT[25]) );
  INV_X1 U21 ( .A(S_IN[25]), .ZN(n8) );
  NAND3_X1 U22 ( .A1(n7), .A2(n6), .A3(\S_IN[15] ), .ZN(n4) );
  NAND2_X1 U23 ( .A1(n4), .A2(n5), .ZN(\S_OUT[26] ) );
  INV_X1 U24 ( .A(EXT_FOR_J), .ZN(n7) );
  INV_X1 U26 ( .A(EXT_UNSIGNED), .ZN(n6) );
endmodule


module register_file_NBIT32_row32 ( CLK, RESET, ENABLE, RD1, RD2, WR, ADD_WR, 
        ADD_RD1, ADD_RD2, DATAIN, OUT1, OUT2 );
  input [4:0] ADD_WR;
  input [4:0] ADD_RD1;
  input [4:0] ADD_RD2;
  input [31:0] DATAIN;
  output [31:0] OUT1;
  output [31:0] OUT2;
  input CLK, RESET, ENABLE, RD1, RD2, WR;
  wire   \REGISTERS[0][31] , \REGISTERS[0][30] , \REGISTERS[0][29] ,
         \REGISTERS[0][28] , \REGISTERS[0][27] , \REGISTERS[0][26] ,
         \REGISTERS[0][25] , \REGISTERS[0][24] , \REGISTERS[0][23] ,
         \REGISTERS[0][22] , \REGISTERS[0][21] , \REGISTERS[0][20] ,
         \REGISTERS[0][19] , \REGISTERS[0][18] , \REGISTERS[0][17] ,
         \REGISTERS[0][16] , \REGISTERS[0][15] , \REGISTERS[0][14] ,
         \REGISTERS[0][13] , \REGISTERS[0][12] , \REGISTERS[0][11] ,
         \REGISTERS[0][10] , \REGISTERS[0][9] , \REGISTERS[0][8] ,
         \REGISTERS[0][7] , \REGISTERS[0][6] , \REGISTERS[0][5] ,
         \REGISTERS[0][4] , \REGISTERS[0][3] , \REGISTERS[0][2] ,
         \REGISTERS[0][1] , \REGISTERS[0][0] , \REGISTERS[1][31] ,
         \REGISTERS[1][30] , \REGISTERS[1][29] , \REGISTERS[1][28] ,
         \REGISTERS[1][27] , \REGISTERS[1][26] , \REGISTERS[1][25] ,
         \REGISTERS[1][24] , \REGISTERS[1][23] , \REGISTERS[1][22] ,
         \REGISTERS[1][21] , \REGISTERS[1][20] , \REGISTERS[1][19] ,
         \REGISTERS[1][18] , \REGISTERS[1][17] , \REGISTERS[1][16] ,
         \REGISTERS[1][15] , \REGISTERS[1][14] , \REGISTERS[1][13] ,
         \REGISTERS[1][12] , \REGISTERS[1][11] , \REGISTERS[1][10] ,
         \REGISTERS[1][9] , \REGISTERS[1][8] , \REGISTERS[1][7] ,
         \REGISTERS[1][6] , \REGISTERS[1][5] , \REGISTERS[1][4] ,
         \REGISTERS[1][3] , \REGISTERS[1][2] , \REGISTERS[1][1] ,
         \REGISTERS[1][0] , \REGISTERS[2][31] , \REGISTERS[2][30] ,
         \REGISTERS[2][29] , \REGISTERS[2][28] , \REGISTERS[2][27] ,
         \REGISTERS[2][26] , \REGISTERS[2][25] , \REGISTERS[2][24] ,
         \REGISTERS[2][23] , \REGISTERS[2][22] , \REGISTERS[2][21] ,
         \REGISTERS[2][20] , \REGISTERS[2][19] , \REGISTERS[2][18] ,
         \REGISTERS[2][17] , \REGISTERS[2][16] , \REGISTERS[2][15] ,
         \REGISTERS[2][14] , \REGISTERS[2][13] , \REGISTERS[2][12] ,
         \REGISTERS[2][11] , \REGISTERS[2][10] , \REGISTERS[2][9] ,
         \REGISTERS[2][8] , \REGISTERS[2][7] , \REGISTERS[2][6] ,
         \REGISTERS[2][5] , \REGISTERS[2][4] , \REGISTERS[2][3] ,
         \REGISTERS[2][2] , \REGISTERS[2][1] , \REGISTERS[2][0] ,
         \REGISTERS[3][31] , \REGISTERS[3][30] , \REGISTERS[3][29] ,
         \REGISTERS[3][28] , \REGISTERS[3][27] , \REGISTERS[3][26] ,
         \REGISTERS[3][25] , \REGISTERS[3][24] , \REGISTERS[3][23] ,
         \REGISTERS[3][22] , \REGISTERS[3][21] , \REGISTERS[3][20] ,
         \REGISTERS[3][19] , \REGISTERS[3][18] , \REGISTERS[3][17] ,
         \REGISTERS[3][16] , \REGISTERS[3][15] , \REGISTERS[3][14] ,
         \REGISTERS[3][13] , \REGISTERS[3][12] , \REGISTERS[3][11] ,
         \REGISTERS[3][10] , \REGISTERS[3][9] , \REGISTERS[3][8] ,
         \REGISTERS[3][7] , \REGISTERS[3][6] , \REGISTERS[3][5] ,
         \REGISTERS[3][4] , \REGISTERS[3][3] , \REGISTERS[3][2] ,
         \REGISTERS[3][1] , \REGISTERS[3][0] , \REGISTERS[4][31] ,
         \REGISTERS[4][30] , \REGISTERS[4][29] , \REGISTERS[4][28] ,
         \REGISTERS[4][27] , \REGISTERS[4][26] , \REGISTERS[4][25] ,
         \REGISTERS[4][24] , \REGISTERS[4][23] , \REGISTERS[4][22] ,
         \REGISTERS[4][21] , \REGISTERS[4][20] , \REGISTERS[4][19] ,
         \REGISTERS[4][18] , \REGISTERS[4][17] , \REGISTERS[4][16] ,
         \REGISTERS[4][15] , \REGISTERS[4][14] , \REGISTERS[4][13] ,
         \REGISTERS[4][12] , \REGISTERS[4][11] , \REGISTERS[4][10] ,
         \REGISTERS[4][9] , \REGISTERS[4][8] , \REGISTERS[4][7] ,
         \REGISTERS[4][6] , \REGISTERS[4][5] , \REGISTERS[4][4] ,
         \REGISTERS[4][3] , \REGISTERS[4][2] , \REGISTERS[4][1] ,
         \REGISTERS[4][0] , \REGISTERS[5][31] , \REGISTERS[5][30] ,
         \REGISTERS[5][29] , \REGISTERS[5][28] , \REGISTERS[5][27] ,
         \REGISTERS[5][26] , \REGISTERS[5][25] , \REGISTERS[5][24] ,
         \REGISTERS[5][23] , \REGISTERS[5][22] , \REGISTERS[5][21] ,
         \REGISTERS[5][20] , \REGISTERS[5][19] , \REGISTERS[5][18] ,
         \REGISTERS[5][17] , \REGISTERS[5][16] , \REGISTERS[5][15] ,
         \REGISTERS[5][14] , \REGISTERS[5][13] , \REGISTERS[5][12] ,
         \REGISTERS[5][11] , \REGISTERS[5][10] , \REGISTERS[5][9] ,
         \REGISTERS[5][8] , \REGISTERS[5][7] , \REGISTERS[5][6] ,
         \REGISTERS[5][5] , \REGISTERS[5][4] , \REGISTERS[5][3] ,
         \REGISTERS[5][2] , \REGISTERS[5][1] , \REGISTERS[5][0] ,
         \REGISTERS[6][31] , \REGISTERS[6][30] , \REGISTERS[6][29] ,
         \REGISTERS[6][28] , \REGISTERS[6][27] , \REGISTERS[6][26] ,
         \REGISTERS[6][25] , \REGISTERS[6][24] , \REGISTERS[6][23] ,
         \REGISTERS[6][22] , \REGISTERS[6][21] , \REGISTERS[6][20] ,
         \REGISTERS[6][19] , \REGISTERS[6][18] , \REGISTERS[6][17] ,
         \REGISTERS[6][16] , \REGISTERS[6][15] , \REGISTERS[6][14] ,
         \REGISTERS[6][13] , \REGISTERS[6][12] , \REGISTERS[6][11] ,
         \REGISTERS[6][10] , \REGISTERS[6][9] , \REGISTERS[6][8] ,
         \REGISTERS[6][7] , \REGISTERS[6][6] , \REGISTERS[6][5] ,
         \REGISTERS[6][4] , \REGISTERS[6][3] , \REGISTERS[6][2] ,
         \REGISTERS[6][1] , \REGISTERS[6][0] , \REGISTERS[7][31] ,
         \REGISTERS[7][30] , \REGISTERS[7][29] , \REGISTERS[7][28] ,
         \REGISTERS[7][27] , \REGISTERS[7][26] , \REGISTERS[7][25] ,
         \REGISTERS[7][24] , \REGISTERS[7][23] , \REGISTERS[7][22] ,
         \REGISTERS[7][21] , \REGISTERS[7][20] , \REGISTERS[7][19] ,
         \REGISTERS[7][18] , \REGISTERS[7][17] , \REGISTERS[7][16] ,
         \REGISTERS[7][15] , \REGISTERS[7][14] , \REGISTERS[7][13] ,
         \REGISTERS[7][12] , \REGISTERS[7][11] , \REGISTERS[7][10] ,
         \REGISTERS[7][9] , \REGISTERS[7][8] , \REGISTERS[7][7] ,
         \REGISTERS[7][6] , \REGISTERS[7][5] , \REGISTERS[7][4] ,
         \REGISTERS[7][3] , \REGISTERS[7][2] , \REGISTERS[7][1] ,
         \REGISTERS[7][0] , \REGISTERS[8][31] , \REGISTERS[8][30] ,
         \REGISTERS[8][29] , \REGISTERS[8][28] , \REGISTERS[8][27] ,
         \REGISTERS[8][26] , \REGISTERS[8][25] , \REGISTERS[8][24] ,
         \REGISTERS[8][23] , \REGISTERS[8][22] , \REGISTERS[8][21] ,
         \REGISTERS[8][20] , \REGISTERS[8][19] , \REGISTERS[8][18] ,
         \REGISTERS[8][17] , \REGISTERS[8][16] , \REGISTERS[8][15] ,
         \REGISTERS[8][14] , \REGISTERS[8][13] , \REGISTERS[8][12] ,
         \REGISTERS[8][11] , \REGISTERS[8][10] , \REGISTERS[8][9] ,
         \REGISTERS[8][8] , \REGISTERS[8][7] , \REGISTERS[8][6] ,
         \REGISTERS[8][5] , \REGISTERS[8][4] , \REGISTERS[8][3] ,
         \REGISTERS[8][2] , \REGISTERS[8][1] , \REGISTERS[8][0] ,
         \REGISTERS[9][31] , \REGISTERS[9][30] , \REGISTERS[9][29] ,
         \REGISTERS[9][28] , \REGISTERS[9][27] , \REGISTERS[9][26] ,
         \REGISTERS[9][25] , \REGISTERS[9][24] , \REGISTERS[9][23] ,
         \REGISTERS[9][22] , \REGISTERS[9][21] , \REGISTERS[9][20] ,
         \REGISTERS[9][19] , \REGISTERS[9][18] , \REGISTERS[9][17] ,
         \REGISTERS[9][16] , \REGISTERS[9][15] , \REGISTERS[9][14] ,
         \REGISTERS[9][13] , \REGISTERS[9][12] , \REGISTERS[9][11] ,
         \REGISTERS[9][10] , \REGISTERS[9][9] , \REGISTERS[9][8] ,
         \REGISTERS[9][7] , \REGISTERS[9][6] , \REGISTERS[9][5] ,
         \REGISTERS[9][4] , \REGISTERS[9][3] , \REGISTERS[9][2] ,
         \REGISTERS[9][1] , \REGISTERS[9][0] , \REGISTERS[10][31] ,
         \REGISTERS[10][30] , \REGISTERS[10][29] , \REGISTERS[10][28] ,
         \REGISTERS[10][27] , \REGISTERS[10][26] , \REGISTERS[10][25] ,
         \REGISTERS[10][24] , \REGISTERS[10][23] , \REGISTERS[10][22] ,
         \REGISTERS[10][21] , \REGISTERS[10][20] , \REGISTERS[10][19] ,
         \REGISTERS[10][18] , \REGISTERS[10][17] , \REGISTERS[10][16] ,
         \REGISTERS[10][15] , \REGISTERS[10][14] , \REGISTERS[10][13] ,
         \REGISTERS[10][12] , \REGISTERS[10][11] , \REGISTERS[10][10] ,
         \REGISTERS[10][9] , \REGISTERS[10][8] , \REGISTERS[10][7] ,
         \REGISTERS[10][6] , \REGISTERS[10][5] , \REGISTERS[10][4] ,
         \REGISTERS[10][3] , \REGISTERS[10][2] , \REGISTERS[10][1] ,
         \REGISTERS[10][0] , \REGISTERS[11][31] , \REGISTERS[11][30] ,
         \REGISTERS[11][29] , \REGISTERS[11][28] , \REGISTERS[11][27] ,
         \REGISTERS[11][26] , \REGISTERS[11][25] , \REGISTERS[11][24] ,
         \REGISTERS[11][23] , \REGISTERS[11][22] , \REGISTERS[11][21] ,
         \REGISTERS[11][20] , \REGISTERS[11][19] , \REGISTERS[11][18] ,
         \REGISTERS[11][17] , \REGISTERS[11][16] , \REGISTERS[11][15] ,
         \REGISTERS[11][14] , \REGISTERS[11][13] , \REGISTERS[11][12] ,
         \REGISTERS[11][11] , \REGISTERS[11][10] , \REGISTERS[11][9] ,
         \REGISTERS[11][8] , \REGISTERS[11][7] , \REGISTERS[11][6] ,
         \REGISTERS[11][5] , \REGISTERS[11][4] , \REGISTERS[11][3] ,
         \REGISTERS[11][2] , \REGISTERS[11][1] , \REGISTERS[11][0] ,
         \REGISTERS[12][31] , \REGISTERS[12][30] , \REGISTERS[12][29] ,
         \REGISTERS[12][28] , \REGISTERS[12][27] , \REGISTERS[12][26] ,
         \REGISTERS[12][25] , \REGISTERS[12][24] , \REGISTERS[12][23] ,
         \REGISTERS[12][22] , \REGISTERS[12][21] , \REGISTERS[12][20] ,
         \REGISTERS[12][19] , \REGISTERS[12][18] , \REGISTERS[12][17] ,
         \REGISTERS[12][16] , \REGISTERS[12][15] , \REGISTERS[12][14] ,
         \REGISTERS[12][13] , \REGISTERS[12][12] , \REGISTERS[12][11] ,
         \REGISTERS[12][10] , \REGISTERS[12][9] , \REGISTERS[12][8] ,
         \REGISTERS[12][7] , \REGISTERS[12][6] , \REGISTERS[12][5] ,
         \REGISTERS[12][4] , \REGISTERS[12][3] , \REGISTERS[12][2] ,
         \REGISTERS[12][1] , \REGISTERS[12][0] , \REGISTERS[13][31] ,
         \REGISTERS[13][30] , \REGISTERS[13][29] , \REGISTERS[13][28] ,
         \REGISTERS[13][27] , \REGISTERS[13][26] , \REGISTERS[13][25] ,
         \REGISTERS[13][24] , \REGISTERS[13][23] , \REGISTERS[13][22] ,
         \REGISTERS[13][21] , \REGISTERS[13][20] , \REGISTERS[13][19] ,
         \REGISTERS[13][18] , \REGISTERS[13][17] , \REGISTERS[13][16] ,
         \REGISTERS[13][15] , \REGISTERS[13][14] , \REGISTERS[13][13] ,
         \REGISTERS[13][12] , \REGISTERS[13][11] , \REGISTERS[13][10] ,
         \REGISTERS[13][9] , \REGISTERS[13][8] , \REGISTERS[13][7] ,
         \REGISTERS[13][6] , \REGISTERS[13][5] , \REGISTERS[13][4] ,
         \REGISTERS[13][3] , \REGISTERS[13][2] , \REGISTERS[13][1] ,
         \REGISTERS[13][0] , \REGISTERS[14][31] , \REGISTERS[14][30] ,
         \REGISTERS[14][29] , \REGISTERS[14][28] , \REGISTERS[14][27] ,
         \REGISTERS[14][26] , \REGISTERS[14][25] , \REGISTERS[14][24] ,
         \REGISTERS[14][23] , \REGISTERS[14][22] , \REGISTERS[14][21] ,
         \REGISTERS[14][20] , \REGISTERS[14][19] , \REGISTERS[14][18] ,
         \REGISTERS[14][17] , \REGISTERS[14][16] , \REGISTERS[14][15] ,
         \REGISTERS[14][14] , \REGISTERS[14][13] , \REGISTERS[14][12] ,
         \REGISTERS[14][11] , \REGISTERS[14][10] , \REGISTERS[14][9] ,
         \REGISTERS[14][8] , \REGISTERS[14][7] , \REGISTERS[14][6] ,
         \REGISTERS[14][5] , \REGISTERS[14][4] , \REGISTERS[14][3] ,
         \REGISTERS[14][2] , \REGISTERS[14][1] , \REGISTERS[14][0] ,
         \REGISTERS[15][31] , \REGISTERS[15][30] , \REGISTERS[15][29] ,
         \REGISTERS[15][28] , \REGISTERS[15][27] , \REGISTERS[15][26] ,
         \REGISTERS[15][25] , \REGISTERS[15][24] , \REGISTERS[15][23] ,
         \REGISTERS[15][22] , \REGISTERS[15][21] , \REGISTERS[15][20] ,
         \REGISTERS[15][19] , \REGISTERS[15][18] , \REGISTERS[15][17] ,
         \REGISTERS[15][16] , \REGISTERS[15][15] , \REGISTERS[15][14] ,
         \REGISTERS[15][13] , \REGISTERS[15][12] , \REGISTERS[15][11] ,
         \REGISTERS[15][10] , \REGISTERS[15][9] , \REGISTERS[15][8] ,
         \REGISTERS[15][7] , \REGISTERS[15][6] , \REGISTERS[15][5] ,
         \REGISTERS[15][4] , \REGISTERS[15][3] , \REGISTERS[15][2] ,
         \REGISTERS[15][1] , \REGISTERS[15][0] , \REGISTERS[16][31] ,
         \REGISTERS[16][30] , \REGISTERS[16][29] , \REGISTERS[16][28] ,
         \REGISTERS[16][27] , \REGISTERS[16][26] , \REGISTERS[16][25] ,
         \REGISTERS[16][24] , \REGISTERS[16][23] , \REGISTERS[16][22] ,
         \REGISTERS[16][21] , \REGISTERS[16][20] , \REGISTERS[16][19] ,
         \REGISTERS[16][18] , \REGISTERS[16][17] , \REGISTERS[16][16] ,
         \REGISTERS[16][15] , \REGISTERS[16][14] , \REGISTERS[16][13] ,
         \REGISTERS[16][12] , \REGISTERS[16][11] , \REGISTERS[16][10] ,
         \REGISTERS[16][9] , \REGISTERS[16][8] , \REGISTERS[16][7] ,
         \REGISTERS[16][6] , \REGISTERS[16][5] , \REGISTERS[16][4] ,
         \REGISTERS[16][3] , \REGISTERS[16][2] , \REGISTERS[16][1] ,
         \REGISTERS[16][0] , \REGISTERS[17][31] , \REGISTERS[17][30] ,
         \REGISTERS[17][29] , \REGISTERS[17][28] , \REGISTERS[17][27] ,
         \REGISTERS[17][26] , \REGISTERS[17][25] , \REGISTERS[17][24] ,
         \REGISTERS[17][23] , \REGISTERS[17][22] , \REGISTERS[17][21] ,
         \REGISTERS[17][20] , \REGISTERS[17][19] , \REGISTERS[17][18] ,
         \REGISTERS[17][17] , \REGISTERS[17][16] , \REGISTERS[17][15] ,
         \REGISTERS[17][14] , \REGISTERS[17][13] , \REGISTERS[17][12] ,
         \REGISTERS[17][11] , \REGISTERS[17][10] , \REGISTERS[17][9] ,
         \REGISTERS[17][8] , \REGISTERS[17][7] , \REGISTERS[17][6] ,
         \REGISTERS[17][5] , \REGISTERS[17][4] , \REGISTERS[17][3] ,
         \REGISTERS[17][2] , \REGISTERS[17][1] , \REGISTERS[17][0] ,
         \REGISTERS[18][31] , \REGISTERS[18][30] , \REGISTERS[18][29] ,
         \REGISTERS[18][28] , \REGISTERS[18][27] , \REGISTERS[18][26] ,
         \REGISTERS[18][25] , \REGISTERS[18][24] , \REGISTERS[18][23] ,
         \REGISTERS[18][22] , \REGISTERS[18][21] , \REGISTERS[18][20] ,
         \REGISTERS[18][19] , \REGISTERS[18][18] , \REGISTERS[18][17] ,
         \REGISTERS[18][16] , \REGISTERS[18][15] , \REGISTERS[18][14] ,
         \REGISTERS[18][13] , \REGISTERS[18][12] , \REGISTERS[18][11] ,
         \REGISTERS[18][10] , \REGISTERS[18][9] , \REGISTERS[18][8] ,
         \REGISTERS[18][7] , \REGISTERS[18][6] , \REGISTERS[18][5] ,
         \REGISTERS[18][4] , \REGISTERS[18][3] , \REGISTERS[18][2] ,
         \REGISTERS[18][1] , \REGISTERS[18][0] , \REGISTERS[19][31] ,
         \REGISTERS[19][30] , \REGISTERS[19][29] , \REGISTERS[19][28] ,
         \REGISTERS[19][27] , \REGISTERS[19][26] , \REGISTERS[19][25] ,
         \REGISTERS[19][24] , \REGISTERS[19][23] , \REGISTERS[19][22] ,
         \REGISTERS[19][21] , \REGISTERS[19][20] , \REGISTERS[19][19] ,
         \REGISTERS[19][18] , \REGISTERS[19][17] , \REGISTERS[19][16] ,
         \REGISTERS[19][15] , \REGISTERS[19][14] , \REGISTERS[19][13] ,
         \REGISTERS[19][12] , \REGISTERS[19][11] , \REGISTERS[19][10] ,
         \REGISTERS[19][9] , \REGISTERS[19][8] , \REGISTERS[19][7] ,
         \REGISTERS[19][6] , \REGISTERS[19][5] , \REGISTERS[19][4] ,
         \REGISTERS[19][3] , \REGISTERS[19][2] , \REGISTERS[19][1] ,
         \REGISTERS[19][0] , \REGISTERS[20][31] , \REGISTERS[20][30] ,
         \REGISTERS[20][29] , \REGISTERS[20][28] , \REGISTERS[20][27] ,
         \REGISTERS[20][26] , \REGISTERS[20][25] , \REGISTERS[20][24] ,
         \REGISTERS[20][23] , \REGISTERS[20][22] , \REGISTERS[20][21] ,
         \REGISTERS[20][20] , \REGISTERS[20][19] , \REGISTERS[20][18] ,
         \REGISTERS[20][17] , \REGISTERS[20][16] , \REGISTERS[20][15] ,
         \REGISTERS[20][14] , \REGISTERS[20][13] , \REGISTERS[20][12] ,
         \REGISTERS[20][11] , \REGISTERS[20][10] , \REGISTERS[20][9] ,
         \REGISTERS[20][8] , \REGISTERS[20][7] , \REGISTERS[20][6] ,
         \REGISTERS[20][5] , \REGISTERS[20][4] , \REGISTERS[20][3] ,
         \REGISTERS[20][2] , \REGISTERS[20][1] , \REGISTERS[20][0] ,
         \REGISTERS[21][31] , \REGISTERS[21][30] , \REGISTERS[21][29] ,
         \REGISTERS[21][28] , \REGISTERS[21][27] , \REGISTERS[21][26] ,
         \REGISTERS[21][25] , \REGISTERS[21][24] , \REGISTERS[21][23] ,
         \REGISTERS[21][22] , \REGISTERS[21][21] , \REGISTERS[21][20] ,
         \REGISTERS[21][19] , \REGISTERS[21][18] , \REGISTERS[21][17] ,
         \REGISTERS[21][16] , \REGISTERS[21][15] , \REGISTERS[21][14] ,
         \REGISTERS[21][13] , \REGISTERS[21][12] , \REGISTERS[21][11] ,
         \REGISTERS[21][10] , \REGISTERS[21][9] , \REGISTERS[21][8] ,
         \REGISTERS[21][7] , \REGISTERS[21][6] , \REGISTERS[21][5] ,
         \REGISTERS[21][4] , \REGISTERS[21][3] , \REGISTERS[21][2] ,
         \REGISTERS[21][1] , \REGISTERS[21][0] , \REGISTERS[22][31] ,
         \REGISTERS[22][30] , \REGISTERS[22][29] , \REGISTERS[22][28] ,
         \REGISTERS[22][27] , \REGISTERS[22][26] , \REGISTERS[22][25] ,
         \REGISTERS[22][24] , \REGISTERS[22][23] , \REGISTERS[22][22] ,
         \REGISTERS[22][21] , \REGISTERS[22][20] , \REGISTERS[22][19] ,
         \REGISTERS[22][18] , \REGISTERS[22][17] , \REGISTERS[22][16] ,
         \REGISTERS[22][15] , \REGISTERS[22][14] , \REGISTERS[22][13] ,
         \REGISTERS[22][12] , \REGISTERS[22][11] , \REGISTERS[22][10] ,
         \REGISTERS[22][9] , \REGISTERS[22][8] , \REGISTERS[22][7] ,
         \REGISTERS[22][6] , \REGISTERS[22][5] , \REGISTERS[22][4] ,
         \REGISTERS[22][3] , \REGISTERS[22][2] , \REGISTERS[22][1] ,
         \REGISTERS[22][0] , \REGISTERS[23][31] , \REGISTERS[23][30] ,
         \REGISTERS[23][29] , \REGISTERS[23][28] , \REGISTERS[23][27] ,
         \REGISTERS[23][26] , \REGISTERS[23][25] , \REGISTERS[23][24] ,
         \REGISTERS[23][23] , \REGISTERS[23][22] , \REGISTERS[23][21] ,
         \REGISTERS[23][20] , \REGISTERS[23][19] , \REGISTERS[23][18] ,
         \REGISTERS[23][17] , \REGISTERS[23][16] , \REGISTERS[23][15] ,
         \REGISTERS[23][14] , \REGISTERS[23][13] , \REGISTERS[23][12] ,
         \REGISTERS[23][11] , \REGISTERS[23][10] , \REGISTERS[23][9] ,
         \REGISTERS[23][8] , \REGISTERS[23][7] , \REGISTERS[23][6] ,
         \REGISTERS[23][5] , \REGISTERS[23][4] , \REGISTERS[23][3] ,
         \REGISTERS[23][2] , \REGISTERS[23][1] , \REGISTERS[23][0] ,
         \REGISTERS[24][31] , \REGISTERS[24][30] , \REGISTERS[24][29] ,
         \REGISTERS[24][28] , \REGISTERS[24][27] , \REGISTERS[24][26] ,
         \REGISTERS[24][25] , \REGISTERS[24][24] , \REGISTERS[24][23] ,
         \REGISTERS[24][22] , \REGISTERS[24][21] , \REGISTERS[24][20] ,
         \REGISTERS[24][19] , \REGISTERS[24][18] , \REGISTERS[24][17] ,
         \REGISTERS[24][16] , \REGISTERS[24][15] , \REGISTERS[24][14] ,
         \REGISTERS[24][13] , \REGISTERS[24][12] , \REGISTERS[24][11] ,
         \REGISTERS[24][10] , \REGISTERS[24][9] , \REGISTERS[24][8] ,
         \REGISTERS[24][7] , \REGISTERS[24][6] , \REGISTERS[24][5] ,
         \REGISTERS[24][4] , \REGISTERS[24][3] , \REGISTERS[24][2] ,
         \REGISTERS[24][1] , \REGISTERS[24][0] , \REGISTERS[25][31] ,
         \REGISTERS[25][30] , \REGISTERS[25][29] , \REGISTERS[25][28] ,
         \REGISTERS[25][27] , \REGISTERS[25][26] , \REGISTERS[25][25] ,
         \REGISTERS[25][24] , \REGISTERS[25][23] , \REGISTERS[25][22] ,
         \REGISTERS[25][21] , \REGISTERS[25][20] , \REGISTERS[25][19] ,
         \REGISTERS[25][18] , \REGISTERS[25][17] , \REGISTERS[25][16] ,
         \REGISTERS[25][15] , \REGISTERS[25][14] , \REGISTERS[25][13] ,
         \REGISTERS[25][12] , \REGISTERS[25][11] , \REGISTERS[25][10] ,
         \REGISTERS[25][9] , \REGISTERS[25][8] , \REGISTERS[25][7] ,
         \REGISTERS[25][6] , \REGISTERS[25][5] , \REGISTERS[25][4] ,
         \REGISTERS[25][3] , \REGISTERS[25][2] , \REGISTERS[25][1] ,
         \REGISTERS[25][0] , \REGISTERS[26][31] , \REGISTERS[26][30] ,
         \REGISTERS[26][29] , \REGISTERS[26][28] , \REGISTERS[26][27] ,
         \REGISTERS[26][26] , \REGISTERS[26][25] , \REGISTERS[26][24] ,
         \REGISTERS[26][23] , \REGISTERS[26][22] , \REGISTERS[26][21] ,
         \REGISTERS[26][20] , \REGISTERS[26][19] , \REGISTERS[26][18] ,
         \REGISTERS[26][17] , \REGISTERS[26][16] , \REGISTERS[26][15] ,
         \REGISTERS[26][14] , \REGISTERS[26][13] , \REGISTERS[26][12] ,
         \REGISTERS[26][11] , \REGISTERS[26][10] , \REGISTERS[26][9] ,
         \REGISTERS[26][8] , \REGISTERS[26][7] , \REGISTERS[26][6] ,
         \REGISTERS[26][5] , \REGISTERS[26][4] , \REGISTERS[26][3] ,
         \REGISTERS[26][2] , \REGISTERS[26][1] , \REGISTERS[26][0] ,
         \REGISTERS[27][31] , \REGISTERS[27][30] , \REGISTERS[27][29] ,
         \REGISTERS[27][28] , \REGISTERS[27][27] , \REGISTERS[27][26] ,
         \REGISTERS[27][25] , \REGISTERS[27][24] , \REGISTERS[27][23] ,
         \REGISTERS[27][22] , \REGISTERS[27][21] , \REGISTERS[27][20] ,
         \REGISTERS[27][19] , \REGISTERS[27][18] , \REGISTERS[27][17] ,
         \REGISTERS[27][16] , \REGISTERS[27][15] , \REGISTERS[27][14] ,
         \REGISTERS[27][13] , \REGISTERS[27][12] , \REGISTERS[27][11] ,
         \REGISTERS[27][10] , \REGISTERS[27][9] , \REGISTERS[27][8] ,
         \REGISTERS[27][7] , \REGISTERS[27][6] , \REGISTERS[27][5] ,
         \REGISTERS[27][4] , \REGISTERS[27][3] , \REGISTERS[27][2] ,
         \REGISTERS[27][1] , \REGISTERS[27][0] , \REGISTERS[28][31] ,
         \REGISTERS[28][30] , \REGISTERS[28][29] , \REGISTERS[28][28] ,
         \REGISTERS[28][27] , \REGISTERS[28][26] , \REGISTERS[28][25] ,
         \REGISTERS[28][24] , \REGISTERS[28][23] , \REGISTERS[28][22] ,
         \REGISTERS[28][21] , \REGISTERS[28][20] , \REGISTERS[28][19] ,
         \REGISTERS[28][18] , \REGISTERS[28][17] , \REGISTERS[28][16] ,
         \REGISTERS[28][15] , \REGISTERS[28][14] , \REGISTERS[28][13] ,
         \REGISTERS[28][12] , \REGISTERS[28][11] , \REGISTERS[28][10] ,
         \REGISTERS[28][9] , \REGISTERS[28][8] , \REGISTERS[28][7] ,
         \REGISTERS[28][6] , \REGISTERS[28][5] , \REGISTERS[28][4] ,
         \REGISTERS[28][3] , \REGISTERS[28][2] , \REGISTERS[28][1] ,
         \REGISTERS[28][0] , \REGISTERS[29][31] , \REGISTERS[29][30] ,
         \REGISTERS[29][29] , \REGISTERS[29][28] , \REGISTERS[29][27] ,
         \REGISTERS[29][26] , \REGISTERS[29][25] , \REGISTERS[29][24] ,
         \REGISTERS[29][23] , \REGISTERS[29][22] , \REGISTERS[29][21] ,
         \REGISTERS[29][20] , \REGISTERS[29][19] , \REGISTERS[29][18] ,
         \REGISTERS[29][17] , \REGISTERS[29][16] , \REGISTERS[29][15] ,
         \REGISTERS[29][14] , \REGISTERS[29][13] , \REGISTERS[29][12] ,
         \REGISTERS[29][11] , \REGISTERS[29][10] , \REGISTERS[29][9] ,
         \REGISTERS[29][8] , \REGISTERS[29][7] , \REGISTERS[29][6] ,
         \REGISTERS[29][5] , \REGISTERS[29][4] , \REGISTERS[29][3] ,
         \REGISTERS[29][2] , \REGISTERS[29][1] , \REGISTERS[29][0] ,
         \REGISTERS[30][31] , \REGISTERS[30][30] , \REGISTERS[30][29] ,
         \REGISTERS[30][28] , \REGISTERS[30][27] , \REGISTERS[30][26] ,
         \REGISTERS[30][25] , \REGISTERS[30][24] , \REGISTERS[30][23] ,
         \REGISTERS[30][22] , \REGISTERS[30][21] , \REGISTERS[30][20] ,
         \REGISTERS[30][19] , \REGISTERS[30][18] , \REGISTERS[30][17] ,
         \REGISTERS[30][16] , \REGISTERS[30][15] , \REGISTERS[30][14] ,
         \REGISTERS[30][13] , \REGISTERS[30][12] , \REGISTERS[30][11] ,
         \REGISTERS[30][10] , \REGISTERS[30][9] , \REGISTERS[30][8] ,
         \REGISTERS[30][7] , \REGISTERS[30][6] , \REGISTERS[30][5] ,
         \REGISTERS[30][4] , \REGISTERS[30][3] , \REGISTERS[30][2] ,
         \REGISTERS[30][1] , \REGISTERS[30][0] , \REGISTERS[31][31] ,
         \REGISTERS[31][30] , \REGISTERS[31][29] , \REGISTERS[31][28] ,
         \REGISTERS[31][27] , \REGISTERS[31][26] , \REGISTERS[31][25] ,
         \REGISTERS[31][24] , \REGISTERS[31][23] , \REGISTERS[31][22] ,
         \REGISTERS[31][21] , \REGISTERS[31][20] , \REGISTERS[31][19] ,
         \REGISTERS[31][18] , \REGISTERS[31][17] , \REGISTERS[31][16] ,
         \REGISTERS[31][15] , \REGISTERS[31][14] , \REGISTERS[31][13] ,
         \REGISTERS[31][12] , \REGISTERS[31][11] , \REGISTERS[31][10] ,
         \REGISTERS[31][9] , \REGISTERS[31][8] , \REGISTERS[31][7] ,
         \REGISTERS[31][6] , \REGISTERS[31][5] , \REGISTERS[31][4] ,
         \REGISTERS[31][3] , \REGISTERS[31][2] , \REGISTERS[31][1] ,
         \REGISTERS[31][0] , N2419, N2421, N2423, N2425, N2427, N2429, N2431,
         N2433, N2435, N2437, N2439, N2441, N2443, N2445, N2447, N2449, N2451,
         N2453, N2455, N2457, N2459, N2461, N2463, N2465, N2467, N2469, N2471,
         N2473, N2475, N2477, N2479, N2481, N2483, N2485, N2487, N2489, N2491,
         N2493, N2495, N2497, N2499, N2501, N2503, N2505, N2507, N2509, N2511,
         N2513, N2515, N2517, N2519, N2521, N2523, N2525, N2527, N2529, N2531,
         N2533, N2535, N2537, N2539, N2541, N2543, N2545, n4352, n4356, n4360,
         n4364, n4368, n4372, n4376, n4380, n4384, n4388, n4392, n4396, n4400,
         n4404, n4408, n4412, n4416, n4420, n4424, n4428, n4432, n4436, n4440,
         n4444, n4448, n4452, n4456, n4460, n4464, n4468, n4472, n4476, n4480,
         n4484, n4488, n4492, n4496, n4500, n4504, n4508, n4512, n4516, n4520,
         n4524, n4528, n4532, n4536, n4540, n4544, n4548, n4552, n4556, n4560,
         n4564, n4568, n4572, n4576, n4580, n4584, n4588, n4592, n4596, n4600,
         n4604, n4608, n4612, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904,
         n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914,
         n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924,
         n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934,
         n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944,
         n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954,
         n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964,
         n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974,
         n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984,
         n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994,
         n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004,
         n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014,
         n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024,
         n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034,
         n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044,
         n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054,
         n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064,
         n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074,
         n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084,
         n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094,
         n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104,
         n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114,
         n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124,
         n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134,
         n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144,
         n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154,
         n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164,
         n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174,
         n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184,
         n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194,
         n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204,
         n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214,
         n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082;
  tri   RD1;
  tri   RD2;

  DLH_X1 \REGISTERS_reg[0][31]  ( .G(n5071), .D(n5072), .Q(\REGISTERS[0][31] )
         );
  DLH_X1 \REGISTERS_reg[0][30]  ( .G(n5069), .D(n5064), .Q(\REGISTERS[0][30] )
         );
  DLH_X1 \REGISTERS_reg[0][29]  ( .G(n5069), .D(n5060), .Q(\REGISTERS[0][29] )
         );
  DLH_X1 \REGISTERS_reg[0][28]  ( .G(n5069), .D(n5056), .Q(\REGISTERS[0][28] )
         );
  DLH_X1 \REGISTERS_reg[0][27]  ( .G(n5069), .D(n5054), .Q(\REGISTERS[0][27] )
         );
  DLH_X1 \REGISTERS_reg[0][26]  ( .G(n5069), .D(n5048), .Q(\REGISTERS[0][26] )
         );
  DLH_X1 \REGISTERS_reg[0][25]  ( .G(n5068), .D(n5044), .Q(\REGISTERS[0][25] )
         );
  DLH_X1 \REGISTERS_reg[0][24]  ( .G(n5069), .D(n5042), .Q(\REGISTERS[0][24] )
         );
  DLH_X1 \REGISTERS_reg[0][23]  ( .G(n5069), .D(n5038), .Q(\REGISTERS[0][23] )
         );
  DLH_X1 \REGISTERS_reg[0][22]  ( .G(n5068), .D(n5032), .Q(\REGISTERS[0][22] )
         );
  DLH_X1 \REGISTERS_reg[0][21]  ( .G(n5068), .D(n5031), .Q(\REGISTERS[0][21] )
         );
  DLH_X1 \REGISTERS_reg[0][20]  ( .G(n5068), .D(n5024), .Q(\REGISTERS[0][20] )
         );
  DLH_X1 \REGISTERS_reg[0][19]  ( .G(n5068), .D(n5022), .Q(\REGISTERS[0][19] )
         );
  DLH_X1 \REGISTERS_reg[0][18]  ( .G(n5070), .D(n5019), .Q(\REGISTERS[0][18] )
         );
  DLH_X1 \REGISTERS_reg[0][17]  ( .G(n5070), .D(n5015), .Q(\REGISTERS[0][17] )
         );
  DLH_X1 \REGISTERS_reg[0][16]  ( .G(n5068), .D(n5011), .Q(\REGISTERS[0][16] )
         );
  DLH_X1 \REGISTERS_reg[0][15]  ( .G(n5070), .D(n5005), .Q(\REGISTERS[0][15] )
         );
  DLH_X1 \REGISTERS_reg[0][14]  ( .G(n5070), .D(n5003), .Q(\REGISTERS[0][14] )
         );
  DLH_X1 \REGISTERS_reg[0][13]  ( .G(n5070), .D(n4998), .Q(\REGISTERS[0][13] )
         );
  DLH_X1 \REGISTERS_reg[0][12]  ( .G(n5068), .D(n4995), .Q(\REGISTERS[0][12] )
         );
  DLH_X1 \REGISTERS_reg[0][11]  ( .G(n5070), .D(n4990), .Q(\REGISTERS[0][11] )
         );
  DLH_X1 \REGISTERS_reg[0][10]  ( .G(n5070), .D(n4987), .Q(\REGISTERS[0][10] )
         );
  DLH_X1 \REGISTERS_reg[0][9]  ( .G(n5069), .D(n4983), .Q(\REGISTERS[0][9] )
         );
  DLH_X1 \REGISTERS_reg[0][8]  ( .G(n5069), .D(n4979), .Q(\REGISTERS[0][8] )
         );
  DLH_X1 \REGISTERS_reg[0][7]  ( .G(n5069), .D(n4972), .Q(\REGISTERS[0][7] )
         );
  DLH_X1 \REGISTERS_reg[0][6]  ( .G(n5068), .D(n4971), .Q(\REGISTERS[0][6] )
         );
  DLH_X1 \REGISTERS_reg[0][5]  ( .G(n5068), .D(n4967), .Q(\REGISTERS[0][5] )
         );
  DLH_X1 \REGISTERS_reg[0][4]  ( .G(n5068), .D(n4960), .Q(\REGISTERS[0][4] )
         );
  DLH_X1 \REGISTERS_reg[0][3]  ( .G(n5070), .D(n4959), .Q(\REGISTERS[0][3] )
         );
  DLH_X1 \REGISTERS_reg[0][2]  ( .G(n5070), .D(n4955), .Q(\REGISTERS[0][2] )
         );
  DLH_X1 \REGISTERS_reg[0][1]  ( .G(n5070), .D(n4950), .Q(\REGISTERS[0][1] )
         );
  DLH_X1 \REGISTERS_reg[0][0]  ( .G(n5071), .D(n4946), .Q(\REGISTERS[0][0] )
         );
  DLH_X1 \REGISTERS_reg[1][31]  ( .G(n4943), .D(n5072), .Q(\REGISTERS[1][31] )
         );
  DLH_X1 \REGISTERS_reg[1][30]  ( .G(n4943), .D(n5064), .Q(\REGISTERS[1][30] )
         );
  DLH_X1 \REGISTERS_reg[1][29]  ( .G(n4941), .D(n5060), .Q(\REGISTERS[1][29] )
         );
  DLH_X1 \REGISTERS_reg[1][28]  ( .G(n4941), .D(n5056), .Q(\REGISTERS[1][28] )
         );
  DLH_X1 \REGISTERS_reg[1][27]  ( .G(n4941), .D(n5052), .Q(\REGISTERS[1][27] )
         );
  DLH_X1 \REGISTERS_reg[1][26]  ( .G(n4941), .D(n5048), .Q(\REGISTERS[1][26] )
         );
  DLH_X1 \REGISTERS_reg[1][25]  ( .G(n4941), .D(n5044), .Q(\REGISTERS[1][25] )
         );
  DLH_X1 \REGISTERS_reg[1][24]  ( .G(n4941), .D(n5040), .Q(\REGISTERS[1][24] )
         );
  DLH_X1 \REGISTERS_reg[1][23]  ( .G(n4941), .D(n5036), .Q(\REGISTERS[1][23] )
         );
  DLH_X1 \REGISTERS_reg[1][22]  ( .G(n4941), .D(n5032), .Q(\REGISTERS[1][22] )
         );
  DLH_X1 \REGISTERS_reg[1][21]  ( .G(n4941), .D(n5031), .Q(\REGISTERS[1][21] )
         );
  DLH_X1 \REGISTERS_reg[1][20]  ( .G(n4941), .D(n5024), .Q(\REGISTERS[1][20] )
         );
  DLH_X1 \REGISTERS_reg[1][19]  ( .G(n4940), .D(n5020), .Q(\REGISTERS[1][19] )
         );
  DLH_X1 \REGISTERS_reg[1][18]  ( .G(n4940), .D(n5019), .Q(\REGISTERS[1][18] )
         );
  DLH_X1 \REGISTERS_reg[1][17]  ( .G(n4940), .D(n5013), .Q(\REGISTERS[1][17] )
         );
  DLH_X1 \REGISTERS_reg[1][16]  ( .G(n4940), .D(n5009), .Q(\REGISTERS[1][16] )
         );
  DLH_X1 \REGISTERS_reg[1][15]  ( .G(n4940), .D(n5005), .Q(\REGISTERS[1][15] )
         );
  DLH_X1 \REGISTERS_reg[1][14]  ( .G(n4940), .D(n5003), .Q(\REGISTERS[1][14] )
         );
  DLH_X1 \REGISTERS_reg[1][13]  ( .G(n4940), .D(n4998), .Q(\REGISTERS[1][13] )
         );
  DLH_X1 \REGISTERS_reg[1][12]  ( .G(n4940), .D(n4993), .Q(\REGISTERS[1][12] )
         );
  DLH_X1 \REGISTERS_reg[1][11]  ( .G(n4940), .D(n4988), .Q(\REGISTERS[1][11] )
         );
  DLH_X1 \REGISTERS_reg[1][10]  ( .G(n4940), .D(n4985), .Q(\REGISTERS[1][10] )
         );
  DLH_X1 \REGISTERS_reg[1][9]  ( .G(n4942), .D(n4981), .Q(\REGISTERS[1][9] )
         );
  DLH_X1 \REGISTERS_reg[1][8]  ( .G(n4942), .D(n4977), .Q(\REGISTERS[1][8] )
         );
  DLH_X1 \REGISTERS_reg[1][7]  ( .G(n4942), .D(n4975), .Q(\REGISTERS[1][7] )
         );
  DLH_X1 \REGISTERS_reg[1][6]  ( .G(n4942), .D(n4969), .Q(\REGISTERS[1][6] )
         );
  DLH_X1 \REGISTERS_reg[1][5]  ( .G(n4942), .D(n4965), .Q(\REGISTERS[1][5] )
         );
  DLH_X1 \REGISTERS_reg[1][4]  ( .G(n4942), .D(n4960), .Q(\REGISTERS[1][4] )
         );
  DLH_X1 \REGISTERS_reg[1][3]  ( .G(n4942), .D(n4959), .Q(\REGISTERS[1][3] )
         );
  DLH_X1 \REGISTERS_reg[1][2]  ( .G(n4942), .D(n4955), .Q(\REGISTERS[1][2] )
         );
  DLH_X1 \REGISTERS_reg[1][1]  ( .G(n4942), .D(n4950), .Q(\REGISTERS[1][1] )
         );
  DLH_X1 \REGISTERS_reg[1][0]  ( .G(n4942), .D(n4945), .Q(\REGISTERS[1][0] )
         );
  DLH_X1 \REGISTERS_reg[2][31]  ( .G(n4939), .D(n5073), .Q(\REGISTERS[2][31] )
         );
  DLH_X1 \REGISTERS_reg[2][30]  ( .G(n4939), .D(n5065), .Q(\REGISTERS[2][30] )
         );
  DLH_X1 \REGISTERS_reg[2][29]  ( .G(n4937), .D(n5061), .Q(\REGISTERS[2][29] )
         );
  DLH_X1 \REGISTERS_reg[2][28]  ( .G(n4937), .D(n5056), .Q(\REGISTERS[2][28] )
         );
  DLH_X1 \REGISTERS_reg[2][27]  ( .G(n4937), .D(n5052), .Q(\REGISTERS[2][27] )
         );
  DLH_X1 \REGISTERS_reg[2][26]  ( .G(n4937), .D(n5049), .Q(\REGISTERS[2][26] )
         );
  DLH_X1 \REGISTERS_reg[2][25]  ( .G(n4937), .D(n5044), .Q(\REGISTERS[2][25] )
         );
  DLH_X1 \REGISTERS_reg[2][24]  ( .G(n4937), .D(n5040), .Q(\REGISTERS[2][24] )
         );
  DLH_X1 \REGISTERS_reg[2][23]  ( .G(n4937), .D(n5036), .Q(\REGISTERS[2][23] )
         );
  DLH_X1 \REGISTERS_reg[2][22]  ( .G(n4937), .D(n5032), .Q(\REGISTERS[2][22] )
         );
  DLH_X1 \REGISTERS_reg[2][21]  ( .G(n4937), .D(n5028), .Q(\REGISTERS[2][21] )
         );
  DLH_X1 \REGISTERS_reg[2][20]  ( .G(n4937), .D(n5024), .Q(\REGISTERS[2][20] )
         );
  DLH_X1 \REGISTERS_reg[2][19]  ( .G(n4936), .D(n5022), .Q(\REGISTERS[2][19] )
         );
  DLH_X1 \REGISTERS_reg[2][18]  ( .G(n4936), .D(n5016), .Q(\REGISTERS[2][18] )
         );
  DLH_X1 \REGISTERS_reg[2][17]  ( .G(n4936), .D(n5014), .Q(\REGISTERS[2][17] )
         );
  DLH_X1 \REGISTERS_reg[2][16]  ( .G(n4936), .D(n5008), .Q(\REGISTERS[2][16] )
         );
  DLH_X1 \REGISTERS_reg[2][15]  ( .G(n4936), .D(n5004), .Q(\REGISTERS[2][15] )
         );
  DLH_X1 \REGISTERS_reg[2][14]  ( .G(n4936), .D(n5000), .Q(\REGISTERS[2][14] )
         );
  DLH_X1 \REGISTERS_reg[2][13]  ( .G(n4936), .D(n4996), .Q(\REGISTERS[2][13] )
         );
  DLH_X1 \REGISTERS_reg[2][12]  ( .G(n4936), .D(n4994), .Q(\REGISTERS[2][12] )
         );
  DLH_X1 \REGISTERS_reg[2][11]  ( .G(n4936), .D(n4990), .Q(\REGISTERS[2][11] )
         );
  DLH_X1 \REGISTERS_reg[2][10]  ( .G(n4936), .D(n4984), .Q(\REGISTERS[2][10] )
         );
  DLH_X1 \REGISTERS_reg[2][9]  ( .G(n4938), .D(n4980), .Q(\REGISTERS[2][9] )
         );
  DLH_X1 \REGISTERS_reg[2][8]  ( .G(n4938), .D(n4978), .Q(\REGISTERS[2][8] )
         );
  DLH_X1 \REGISTERS_reg[2][7]  ( .G(n4938), .D(n4974), .Q(\REGISTERS[2][7] )
         );
  DLH_X1 \REGISTERS_reg[2][6]  ( .G(n4938), .D(n4970), .Q(\REGISTERS[2][6] )
         );
  DLH_X1 \REGISTERS_reg[2][5]  ( .G(n4938), .D(n4966), .Q(\REGISTERS[2][5] )
         );
  DLH_X1 \REGISTERS_reg[2][4]  ( .G(n4938), .D(n4961), .Q(\REGISTERS[2][4] )
         );
  DLH_X1 \REGISTERS_reg[2][3]  ( .G(n4938), .D(n4956), .Q(\REGISTERS[2][3] )
         );
  DLH_X1 \REGISTERS_reg[2][2]  ( .G(n4938), .D(n4952), .Q(\REGISTERS[2][2] )
         );
  DLH_X1 \REGISTERS_reg[2][1]  ( .G(n4938), .D(n4948), .Q(\REGISTERS[2][1] )
         );
  DLH_X1 \REGISTERS_reg[2][0]  ( .G(n4938), .D(n4946), .Q(\REGISTERS[2][0] )
         );
  DLH_X1 \REGISTERS_reg[3][31]  ( .G(n4935), .D(n5072), .Q(\REGISTERS[3][31] )
         );
  DLH_X1 \REGISTERS_reg[3][30]  ( .G(n4935), .D(n5065), .Q(\REGISTERS[3][30] )
         );
  DLH_X1 \REGISTERS_reg[3][29]  ( .G(n4933), .D(n5061), .Q(\REGISTERS[3][29] )
         );
  DLH_X1 \REGISTERS_reg[3][28]  ( .G(n4933), .D(n5057), .Q(\REGISTERS[3][28] )
         );
  DLH_X1 \REGISTERS_reg[3][27]  ( .G(n4933), .D(n5052), .Q(\REGISTERS[3][27] )
         );
  DLH_X1 \REGISTERS_reg[3][26]  ( .G(n4933), .D(n5049), .Q(\REGISTERS[3][26] )
         );
  DLH_X1 \REGISTERS_reg[3][25]  ( .G(n4933), .D(n5045), .Q(\REGISTERS[3][25] )
         );
  DLH_X1 \REGISTERS_reg[3][24]  ( .G(n4933), .D(n5040), .Q(\REGISTERS[3][24] )
         );
  DLH_X1 \REGISTERS_reg[3][23]  ( .G(n4933), .D(n5036), .Q(\REGISTERS[3][23] )
         );
  DLH_X1 \REGISTERS_reg[3][22]  ( .G(n4933), .D(n5033), .Q(\REGISTERS[3][22] )
         );
  DLH_X1 \REGISTERS_reg[3][21]  ( .G(n4933), .D(n5029), .Q(\REGISTERS[3][21] )
         );
  DLH_X1 \REGISTERS_reg[3][20]  ( .G(n4933), .D(n5025), .Q(\REGISTERS[3][20] )
         );
  DLH_X1 \REGISTERS_reg[3][19]  ( .G(n4932), .D(n5023), .Q(\REGISTERS[3][19] )
         );
  DLH_X1 \REGISTERS_reg[3][18]  ( .G(n4932), .D(n5017), .Q(\REGISTERS[3][18] )
         );
  DLH_X1 \REGISTERS_reg[3][17]  ( .G(n4932), .D(n5013), .Q(\REGISTERS[3][17] )
         );
  DLH_X1 \REGISTERS_reg[3][16]  ( .G(n4932), .D(n5009), .Q(\REGISTERS[3][16] )
         );
  DLH_X1 \REGISTERS_reg[3][15]  ( .G(n4932), .D(n5006), .Q(\REGISTERS[3][15] )
         );
  DLH_X1 \REGISTERS_reg[3][14]  ( .G(n4932), .D(n5001), .Q(\REGISTERS[3][14] )
         );
  DLH_X1 \REGISTERS_reg[3][13]  ( .G(n4932), .D(n4997), .Q(\REGISTERS[3][13] )
         );
  DLH_X1 \REGISTERS_reg[3][12]  ( .G(n4932), .D(n4993), .Q(\REGISTERS[3][12] )
         );
  DLH_X1 \REGISTERS_reg[3][11]  ( .G(n4932), .D(n4990), .Q(\REGISTERS[3][11] )
         );
  DLH_X1 \REGISTERS_reg[3][10]  ( .G(n4932), .D(n4985), .Q(\REGISTERS[3][10] )
         );
  DLH_X1 \REGISTERS_reg[3][9]  ( .G(n4934), .D(n4981), .Q(\REGISTERS[3][9] )
         );
  DLH_X1 \REGISTERS_reg[3][8]  ( .G(n4934), .D(n4977), .Q(\REGISTERS[3][8] )
         );
  DLH_X1 \REGISTERS_reg[3][7]  ( .G(n4934), .D(n4973), .Q(\REGISTERS[3][7] )
         );
  DLH_X1 \REGISTERS_reg[3][6]  ( .G(n4934), .D(n4969), .Q(\REGISTERS[3][6] )
         );
  DLH_X1 \REGISTERS_reg[3][5]  ( .G(n4934), .D(n4965), .Q(\REGISTERS[3][5] )
         );
  DLH_X1 \REGISTERS_reg[3][4]  ( .G(n4934), .D(n4960), .Q(\REGISTERS[3][4] )
         );
  DLH_X1 \REGISTERS_reg[3][3]  ( .G(n4934), .D(n4957), .Q(\REGISTERS[3][3] )
         );
  DLH_X1 \REGISTERS_reg[3][2]  ( .G(n4934), .D(n4953), .Q(\REGISTERS[3][2] )
         );
  DLH_X1 \REGISTERS_reg[3][1]  ( .G(n4934), .D(n4949), .Q(\REGISTERS[3][1] )
         );
  DLH_X1 \REGISTERS_reg[3][0]  ( .G(n4934), .D(n4945), .Q(\REGISTERS[3][0] )
         );
  DLH_X1 \REGISTERS_reg[4][31]  ( .G(n4931), .D(n5072), .Q(\REGISTERS[4][31] )
         );
  DLH_X1 \REGISTERS_reg[4][30]  ( .G(n4931), .D(n5064), .Q(\REGISTERS[4][30] )
         );
  DLH_X1 \REGISTERS_reg[4][29]  ( .G(n4929), .D(n5060), .Q(\REGISTERS[4][29] )
         );
  DLH_X1 \REGISTERS_reg[4][28]  ( .G(n4929), .D(n5058), .Q(\REGISTERS[4][28] )
         );
  DLH_X1 \REGISTERS_reg[4][27]  ( .G(n4929), .D(n5052), .Q(\REGISTERS[4][27] )
         );
  DLH_X1 \REGISTERS_reg[4][26]  ( .G(n4929), .D(n5048), .Q(\REGISTERS[4][26] )
         );
  DLH_X1 \REGISTERS_reg[4][25]  ( .G(n4929), .D(n5046), .Q(\REGISTERS[4][25] )
         );
  DLH_X1 \REGISTERS_reg[4][24]  ( .G(n4929), .D(n5041), .Q(\REGISTERS[4][24] )
         );
  DLH_X1 \REGISTERS_reg[4][23]  ( .G(n4929), .D(n5036), .Q(\REGISTERS[4][23] )
         );
  DLH_X1 \REGISTERS_reg[4][22]  ( .G(n4929), .D(n5034), .Q(\REGISTERS[4][22] )
         );
  DLH_X1 \REGISTERS_reg[4][21]  ( .G(n4929), .D(n5028), .Q(\REGISTERS[4][21] )
         );
  DLH_X1 \REGISTERS_reg[4][20]  ( .G(n4929), .D(n5026), .Q(\REGISTERS[4][20] )
         );
  DLH_X1 \REGISTERS_reg[4][19]  ( .G(n4928), .D(n5020), .Q(\REGISTERS[4][19] )
         );
  DLH_X1 \REGISTERS_reg[4][18]  ( .G(n4928), .D(n5016), .Q(\REGISTERS[4][18] )
         );
  DLH_X1 \REGISTERS_reg[4][17]  ( .G(n4928), .D(n5012), .Q(\REGISTERS[4][17] )
         );
  DLH_X1 \REGISTERS_reg[4][16]  ( .G(n4928), .D(n5009), .Q(\REGISTERS[4][16] )
         );
  DLH_X1 \REGISTERS_reg[4][15]  ( .G(n4928), .D(n5004), .Q(\REGISTERS[4][15] )
         );
  DLH_X1 \REGISTERS_reg[4][14]  ( .G(n4928), .D(n5000), .Q(\REGISTERS[4][14] )
         );
  DLH_X1 \REGISTERS_reg[4][13]  ( .G(n4928), .D(n4996), .Q(\REGISTERS[4][13] )
         );
  DLH_X1 \REGISTERS_reg[4][12]  ( .G(n4928), .D(n4992), .Q(\REGISTERS[4][12] )
         );
  DLH_X1 \REGISTERS_reg[4][11]  ( .G(n4928), .D(n4988), .Q(\REGISTERS[4][11] )
         );
  DLH_X1 \REGISTERS_reg[4][10]  ( .G(n4928), .D(n4985), .Q(\REGISTERS[4][10] )
         );
  DLH_X1 \REGISTERS_reg[4][9]  ( .G(n4930), .D(n4981), .Q(\REGISTERS[4][9] )
         );
  DLH_X1 \REGISTERS_reg[4][8]  ( .G(n4930), .D(n4976), .Q(\REGISTERS[4][8] )
         );
  DLH_X1 \REGISTERS_reg[4][7]  ( .G(n4930), .D(n4972), .Q(\REGISTERS[4][7] )
         );
  DLH_X1 \REGISTERS_reg[4][6]  ( .G(n4930), .D(n4968), .Q(\REGISTERS[4][6] )
         );
  DLH_X1 \REGISTERS_reg[4][5]  ( .G(n4930), .D(n4964), .Q(\REGISTERS[4][5] )
         );
  DLH_X1 \REGISTERS_reg[4][4]  ( .G(n4930), .D(n4961), .Q(\REGISTERS[4][4] )
         );
  DLH_X1 \REGISTERS_reg[4][3]  ( .G(n4930), .D(n4956), .Q(\REGISTERS[4][3] )
         );
  DLH_X1 \REGISTERS_reg[4][2]  ( .G(n4930), .D(n4952), .Q(\REGISTERS[4][2] )
         );
  DLH_X1 \REGISTERS_reg[4][1]  ( .G(n4930), .D(n4948), .Q(\REGISTERS[4][1] )
         );
  DLH_X1 \REGISTERS_reg[4][0]  ( .G(n4930), .D(n4944), .Q(\REGISTERS[4][0] )
         );
  DLH_X1 \REGISTERS_reg[5][31]  ( .G(n4927), .D(n5072), .Q(\REGISTERS[5][31] )
         );
  DLH_X1 \REGISTERS_reg[5][30]  ( .G(n4927), .D(n5066), .Q(\REGISTERS[5][30] )
         );
  DLH_X1 \REGISTERS_reg[5][29]  ( .G(n4925), .D(n5062), .Q(\REGISTERS[5][29] )
         );
  DLH_X1 \REGISTERS_reg[5][28]  ( .G(n4925), .D(n5058), .Q(\REGISTERS[5][28] )
         );
  DLH_X1 \REGISTERS_reg[5][27]  ( .G(n4925), .D(n5052), .Q(\REGISTERS[5][27] )
         );
  DLH_X1 \REGISTERS_reg[5][26]  ( .G(n4925), .D(n5050), .Q(\REGISTERS[5][26] )
         );
  DLH_X1 \REGISTERS_reg[5][25]  ( .G(n4925), .D(n5046), .Q(\REGISTERS[5][25] )
         );
  DLH_X1 \REGISTERS_reg[5][24]  ( .G(n4925), .D(n5041), .Q(\REGISTERS[5][24] )
         );
  DLH_X1 \REGISTERS_reg[5][23]  ( .G(n4925), .D(n5036), .Q(\REGISTERS[5][23] )
         );
  DLH_X1 \REGISTERS_reg[5][22]  ( .G(n4925), .D(n5034), .Q(\REGISTERS[5][22] )
         );
  DLH_X1 \REGISTERS_reg[5][21]  ( .G(n4925), .D(n5028), .Q(\REGISTERS[5][21] )
         );
  DLH_X1 \REGISTERS_reg[5][20]  ( .G(n4925), .D(n5026), .Q(\REGISTERS[5][20] )
         );
  DLH_X1 \REGISTERS_reg[5][19]  ( .G(n4924), .D(n5021), .Q(\REGISTERS[5][19] )
         );
  DLH_X1 \REGISTERS_reg[5][18]  ( .G(n4924), .D(n5016), .Q(\REGISTERS[5][18] )
         );
  DLH_X1 \REGISTERS_reg[5][17]  ( .G(n4924), .D(n5013), .Q(\REGISTERS[5][17] )
         );
  DLH_X1 \REGISTERS_reg[5][16]  ( .G(n4924), .D(n5009), .Q(\REGISTERS[5][16] )
         );
  DLH_X1 \REGISTERS_reg[5][15]  ( .G(n4924), .D(n5006), .Q(\REGISTERS[5][15] )
         );
  DLH_X1 \REGISTERS_reg[5][14]  ( .G(n4924), .D(n5000), .Q(\REGISTERS[5][14] )
         );
  DLH_X1 \REGISTERS_reg[5][13]  ( .G(n4924), .D(n4996), .Q(\REGISTERS[5][13] )
         );
  DLH_X1 \REGISTERS_reg[5][12]  ( .G(n4924), .D(n4993), .Q(\REGISTERS[5][12] )
         );
  DLH_X1 \REGISTERS_reg[5][11]  ( .G(n4924), .D(n4988), .Q(\REGISTERS[5][11] )
         );
  DLH_X1 \REGISTERS_reg[5][10]  ( .G(n4924), .D(n4985), .Q(\REGISTERS[5][10] )
         );
  DLH_X1 \REGISTERS_reg[5][9]  ( .G(n4926), .D(n4981), .Q(\REGISTERS[5][9] )
         );
  DLH_X1 \REGISTERS_reg[5][8]  ( .G(n4926), .D(n4977), .Q(\REGISTERS[5][8] )
         );
  DLH_X1 \REGISTERS_reg[5][7]  ( .G(n4926), .D(n4973), .Q(\REGISTERS[5][7] )
         );
  DLH_X1 \REGISTERS_reg[5][6]  ( .G(n4926), .D(n4969), .Q(\REGISTERS[5][6] )
         );
  DLH_X1 \REGISTERS_reg[5][5]  ( .G(n4926), .D(n4965), .Q(\REGISTERS[5][5] )
         );
  DLH_X1 \REGISTERS_reg[5][4]  ( .G(n4926), .D(n4961), .Q(\REGISTERS[5][4] )
         );
  DLH_X1 \REGISTERS_reg[5][3]  ( .G(n4926), .D(n4956), .Q(\REGISTERS[5][3] )
         );
  DLH_X1 \REGISTERS_reg[5][2]  ( .G(n4926), .D(n4952), .Q(\REGISTERS[5][2] )
         );
  DLH_X1 \REGISTERS_reg[5][1]  ( .G(n4926), .D(n4948), .Q(\REGISTERS[5][1] )
         );
  DLH_X1 \REGISTERS_reg[5][0]  ( .G(n4926), .D(n4945), .Q(\REGISTERS[5][0] )
         );
  DLH_X1 \REGISTERS_reg[6][31]  ( .G(n4923), .D(n5074), .Q(\REGISTERS[6][31] )
         );
  DLH_X1 \REGISTERS_reg[6][30]  ( .G(n4923), .D(n5066), .Q(\REGISTERS[6][30] )
         );
  DLH_X1 \REGISTERS_reg[6][29]  ( .G(n4921), .D(n5062), .Q(\REGISTERS[6][29] )
         );
  DLH_X1 \REGISTERS_reg[6][28]  ( .G(n4921), .D(n5057), .Q(\REGISTERS[6][28] )
         );
  DLH_X1 \REGISTERS_reg[6][27]  ( .G(n4921), .D(n5054), .Q(\REGISTERS[6][27] )
         );
  DLH_X1 \REGISTERS_reg[6][26]  ( .G(n4921), .D(n5050), .Q(\REGISTERS[6][26] )
         );
  DLH_X1 \REGISTERS_reg[6][25]  ( .G(n4921), .D(n5045), .Q(\REGISTERS[6][25] )
         );
  DLH_X1 \REGISTERS_reg[6][24]  ( .G(n4921), .D(n5042), .Q(\REGISTERS[6][24] )
         );
  DLH_X1 \REGISTERS_reg[6][23]  ( .G(n4921), .D(n5038), .Q(\REGISTERS[6][23] )
         );
  DLH_X1 \REGISTERS_reg[6][22]  ( .G(n4921), .D(n5033), .Q(\REGISTERS[6][22] )
         );
  DLH_X1 \REGISTERS_reg[6][21]  ( .G(n4921), .D(n5029), .Q(\REGISTERS[6][21] )
         );
  DLH_X1 \REGISTERS_reg[6][20]  ( .G(n4921), .D(n5025), .Q(\REGISTERS[6][20] )
         );
  DLH_X1 \REGISTERS_reg[6][19]  ( .G(n4920), .D(n5020), .Q(\REGISTERS[6][19] )
         );
  DLH_X1 \REGISTERS_reg[6][18]  ( .G(n4920), .D(n5017), .Q(\REGISTERS[6][18] )
         );
  DLH_X1 \REGISTERS_reg[6][17]  ( .G(n4920), .D(n5012), .Q(\REGISTERS[6][17] )
         );
  DLH_X1 \REGISTERS_reg[6][16]  ( .G(n4920), .D(n5011), .Q(\REGISTERS[6][16] )
         );
  DLH_X1 \REGISTERS_reg[6][15]  ( .G(n4920), .D(n5006), .Q(\REGISTERS[6][15] )
         );
  DLH_X1 \REGISTERS_reg[6][14]  ( .G(n4920), .D(n5001), .Q(\REGISTERS[6][14] )
         );
  DLH_X1 \REGISTERS_reg[6][13]  ( .G(n4920), .D(n4997), .Q(\REGISTERS[6][13] )
         );
  DLH_X1 \REGISTERS_reg[6][12]  ( .G(n4920), .D(n4992), .Q(\REGISTERS[6][12] )
         );
  DLH_X1 \REGISTERS_reg[6][11]  ( .G(n4920), .D(n4988), .Q(\REGISTERS[6][11] )
         );
  DLH_X1 \REGISTERS_reg[6][10]  ( .G(n4920), .D(n4987), .Q(\REGISTERS[6][10] )
         );
  DLH_X1 \REGISTERS_reg[6][9]  ( .G(n4922), .D(n4983), .Q(\REGISTERS[6][9] )
         );
  DLH_X1 \REGISTERS_reg[6][8]  ( .G(n4922), .D(n4976), .Q(\REGISTERS[6][8] )
         );
  DLH_X1 \REGISTERS_reg[6][7]  ( .G(n4922), .D(n4972), .Q(\REGISTERS[6][7] )
         );
  DLH_X1 \REGISTERS_reg[6][6]  ( .G(n4922), .D(n4968), .Q(\REGISTERS[6][6] )
         );
  DLH_X1 \REGISTERS_reg[6][5]  ( .G(n4922), .D(n4964), .Q(\REGISTERS[6][5] )
         );
  DLH_X1 \REGISTERS_reg[6][4]  ( .G(n4922), .D(n4963), .Q(\REGISTERS[6][4] )
         );
  DLH_X1 \REGISTERS_reg[6][3]  ( .G(n4922), .D(n4957), .Q(\REGISTERS[6][3] )
         );
  DLH_X1 \REGISTERS_reg[6][2]  ( .G(n4922), .D(n4953), .Q(\REGISTERS[6][2] )
         );
  DLH_X1 \REGISTERS_reg[6][1]  ( .G(n4922), .D(n4949), .Q(\REGISTERS[6][1] )
         );
  DLH_X1 \REGISTERS_reg[6][0]  ( .G(n4922), .D(n4944), .Q(\REGISTERS[6][0] )
         );
  DLH_X1 \REGISTERS_reg[7][31]  ( .G(n4919), .D(n5074), .Q(\REGISTERS[7][31] )
         );
  DLH_X1 \REGISTERS_reg[7][30]  ( .G(n4919), .D(n5064), .Q(\REGISTERS[7][30] )
         );
  DLH_X1 \REGISTERS_reg[7][29]  ( .G(n4917), .D(n5060), .Q(\REGISTERS[7][29] )
         );
  DLH_X1 \REGISTERS_reg[7][28]  ( .G(n4917), .D(n5057), .Q(\REGISTERS[7][28] )
         );
  DLH_X1 \REGISTERS_reg[7][27]  ( .G(n4917), .D(n5054), .Q(\REGISTERS[7][27] )
         );
  DLH_X1 \REGISTERS_reg[7][26]  ( .G(n4917), .D(n5048), .Q(\REGISTERS[7][26] )
         );
  DLH_X1 \REGISTERS_reg[7][25]  ( .G(n4917), .D(n5045), .Q(\REGISTERS[7][25] )
         );
  DLH_X1 \REGISTERS_reg[7][24]  ( .G(n4917), .D(n5042), .Q(\REGISTERS[7][24] )
         );
  DLH_X1 \REGISTERS_reg[7][23]  ( .G(n4917), .D(n5038), .Q(\REGISTERS[7][23] )
         );
  DLH_X1 \REGISTERS_reg[7][22]  ( .G(n4917), .D(n5033), .Q(\REGISTERS[7][22] )
         );
  DLH_X1 \REGISTERS_reg[7][21]  ( .G(n4917), .D(n5030), .Q(\REGISTERS[7][21] )
         );
  DLH_X1 \REGISTERS_reg[7][20]  ( .G(n4917), .D(n5025), .Q(\REGISTERS[7][20] )
         );
  DLH_X1 \REGISTERS_reg[7][19]  ( .G(n4916), .D(n5020), .Q(\REGISTERS[7][19] )
         );
  DLH_X1 \REGISTERS_reg[7][18]  ( .G(n4916), .D(n5018), .Q(\REGISTERS[7][18] )
         );
  DLH_X1 \REGISTERS_reg[7][17]  ( .G(n4916), .D(n5014), .Q(\REGISTERS[7][17] )
         );
  DLH_X1 \REGISTERS_reg[7][16]  ( .G(n4916), .D(n5010), .Q(\REGISTERS[7][16] )
         );
  DLH_X1 \REGISTERS_reg[7][15]  ( .G(n4916), .D(n5006), .Q(\REGISTERS[7][15] )
         );
  DLH_X1 \REGISTERS_reg[7][14]  ( .G(n4916), .D(n5002), .Q(\REGISTERS[7][14] )
         );
  DLH_X1 \REGISTERS_reg[7][13]  ( .G(n4916), .D(n4998), .Q(\REGISTERS[7][13] )
         );
  DLH_X1 \REGISTERS_reg[7][12]  ( .G(n4916), .D(n4994), .Q(\REGISTERS[7][12] )
         );
  DLH_X1 \REGISTERS_reg[7][11]  ( .G(n4916), .D(n4988), .Q(\REGISTERS[7][11] )
         );
  DLH_X1 \REGISTERS_reg[7][10]  ( .G(n4916), .D(n4986), .Q(\REGISTERS[7][10] )
         );
  DLH_X1 \REGISTERS_reg[7][9]  ( .G(n4918), .D(n4982), .Q(\REGISTERS[7][9] )
         );
  DLH_X1 \REGISTERS_reg[7][8]  ( .G(n4918), .D(n4978), .Q(\REGISTERS[7][8] )
         );
  DLH_X1 \REGISTERS_reg[7][7]  ( .G(n4918), .D(n4972), .Q(\REGISTERS[7][7] )
         );
  DLH_X1 \REGISTERS_reg[7][6]  ( .G(n4918), .D(n4970), .Q(\REGISTERS[7][6] )
         );
  DLH_X1 \REGISTERS_reg[7][5]  ( .G(n4918), .D(n4966), .Q(\REGISTERS[7][5] )
         );
  DLH_X1 \REGISTERS_reg[7][4]  ( .G(n4918), .D(n4963), .Q(\REGISTERS[7][4] )
         );
  DLH_X1 \REGISTERS_reg[7][3]  ( .G(n4918), .D(n4958), .Q(\REGISTERS[7][3] )
         );
  DLH_X1 \REGISTERS_reg[7][2]  ( .G(n4918), .D(n4954), .Q(\REGISTERS[7][2] )
         );
  DLH_X1 \REGISTERS_reg[7][1]  ( .G(n4918), .D(n4950), .Q(\REGISTERS[7][1] )
         );
  DLH_X1 \REGISTERS_reg[7][0]  ( .G(n4918), .D(n4945), .Q(\REGISTERS[7][0] )
         );
  DLH_X1 \REGISTERS_reg[8][31]  ( .G(n4915), .D(n5074), .Q(\REGISTERS[8][31] )
         );
  DLH_X1 \REGISTERS_reg[8][30]  ( .G(n4915), .D(n5066), .Q(\REGISTERS[8][30] )
         );
  DLH_X1 \REGISTERS_reg[8][29]  ( .G(n4913), .D(n5062), .Q(\REGISTERS[8][29] )
         );
  DLH_X1 \REGISTERS_reg[8][28]  ( .G(n4913), .D(n5058), .Q(\REGISTERS[8][28] )
         );
  DLH_X1 \REGISTERS_reg[8][27]  ( .G(n4913), .D(n5054), .Q(\REGISTERS[8][27] )
         );
  DLH_X1 \REGISTERS_reg[8][26]  ( .G(n4913), .D(n5050), .Q(\REGISTERS[8][26] )
         );
  DLH_X1 \REGISTERS_reg[8][25]  ( .G(n4913), .D(n5046), .Q(\REGISTERS[8][25] )
         );
  DLH_X1 \REGISTERS_reg[8][24]  ( .G(n4913), .D(n5042), .Q(\REGISTERS[8][24] )
         );
  DLH_X1 \REGISTERS_reg[8][23]  ( .G(n4913), .D(n5038), .Q(\REGISTERS[8][23] )
         );
  DLH_X1 \REGISTERS_reg[8][22]  ( .G(n4913), .D(n5034), .Q(\REGISTERS[8][22] )
         );
  DLH_X1 \REGISTERS_reg[8][21]  ( .G(n4913), .D(n5030), .Q(\REGISTERS[8][21] )
         );
  DLH_X1 \REGISTERS_reg[8][20]  ( .G(n4913), .D(n5026), .Q(\REGISTERS[8][20] )
         );
  DLH_X1 \REGISTERS_reg[8][19]  ( .G(n4912), .D(n5022), .Q(\REGISTERS[8][19] )
         );
  DLH_X1 \REGISTERS_reg[8][18]  ( .G(n4912), .D(n5018), .Q(\REGISTERS[8][18] )
         );
  DLH_X1 \REGISTERS_reg[8][17]  ( .G(n4912), .D(n5014), .Q(\REGISTERS[8][17] )
         );
  DLH_X1 \REGISTERS_reg[8][16]  ( .G(n4912), .D(n5010), .Q(\REGISTERS[8][16] )
         );
  DLH_X1 \REGISTERS_reg[8][15]  ( .G(n4912), .D(n5006), .Q(\REGISTERS[8][15] )
         );
  DLH_X1 \REGISTERS_reg[8][14]  ( .G(n4912), .D(n5002), .Q(\REGISTERS[8][14] )
         );
  DLH_X1 \REGISTERS_reg[8][13]  ( .G(n4912), .D(n4998), .Q(\REGISTERS[8][13] )
         );
  DLH_X1 \REGISTERS_reg[8][12]  ( .G(n4912), .D(n4994), .Q(\REGISTERS[8][12] )
         );
  DLH_X1 \REGISTERS_reg[8][11]  ( .G(n4912), .D(n4990), .Q(\REGISTERS[8][11] )
         );
  DLH_X1 \REGISTERS_reg[8][10]  ( .G(n4912), .D(n4986), .Q(\REGISTERS[8][10] )
         );
  DLH_X1 \REGISTERS_reg[8][9]  ( .G(n4914), .D(n4982), .Q(\REGISTERS[8][9] )
         );
  DLH_X1 \REGISTERS_reg[8][8]  ( .G(n4914), .D(n4978), .Q(\REGISTERS[8][8] )
         );
  DLH_X1 \REGISTERS_reg[8][7]  ( .G(n4914), .D(n4974), .Q(\REGISTERS[8][7] )
         );
  DLH_X1 \REGISTERS_reg[8][6]  ( .G(n4914), .D(n4970), .Q(\REGISTERS[8][6] )
         );
  DLH_X1 \REGISTERS_reg[8][5]  ( .G(n4914), .D(n4966), .Q(\REGISTERS[8][5] )
         );
  DLH_X1 \REGISTERS_reg[8][4]  ( .G(n4914), .D(n4962), .Q(\REGISTERS[8][4] )
         );
  DLH_X1 \REGISTERS_reg[8][3]  ( .G(n4914), .D(n4958), .Q(\REGISTERS[8][3] )
         );
  DLH_X1 \REGISTERS_reg[8][2]  ( .G(n4914), .D(n4954), .Q(\REGISTERS[8][2] )
         );
  DLH_X1 \REGISTERS_reg[8][1]  ( .G(n4914), .D(n4950), .Q(\REGISTERS[8][1] )
         );
  DLH_X1 \REGISTERS_reg[8][0]  ( .G(n4914), .D(n4946), .Q(\REGISTERS[8][0] )
         );
  DLH_X1 \REGISTERS_reg[9][31]  ( .G(n4911), .D(n5072), .Q(\REGISTERS[9][31] )
         );
  DLH_X1 \REGISTERS_reg[9][30]  ( .G(n4911), .D(n5065), .Q(\REGISTERS[9][30] )
         );
  DLH_X1 \REGISTERS_reg[9][29]  ( .G(n4909), .D(n5061), .Q(\REGISTERS[9][29] )
         );
  DLH_X1 \REGISTERS_reg[9][28]  ( .G(n4909), .D(n5057), .Q(\REGISTERS[9][28] )
         );
  DLH_X1 \REGISTERS_reg[9][27]  ( .G(n4909), .D(n5053), .Q(\REGISTERS[9][27] )
         );
  DLH_X1 \REGISTERS_reg[9][26]  ( .G(n4909), .D(n5049), .Q(\REGISTERS[9][26] )
         );
  DLH_X1 \REGISTERS_reg[9][25]  ( .G(n4909), .D(n5045), .Q(\REGISTERS[9][25] )
         );
  DLH_X1 \REGISTERS_reg[9][24]  ( .G(n4909), .D(n5040), .Q(\REGISTERS[9][24] )
         );
  DLH_X1 \REGISTERS_reg[9][23]  ( .G(n4909), .D(n5037), .Q(\REGISTERS[9][23] )
         );
  DLH_X1 \REGISTERS_reg[9][22]  ( .G(n4909), .D(n5033), .Q(\REGISTERS[9][22] )
         );
  DLH_X1 \REGISTERS_reg[9][21]  ( .G(n4909), .D(n5029), .Q(\REGISTERS[9][21] )
         );
  DLH_X1 \REGISTERS_reg[9][20]  ( .G(n4909), .D(n5025), .Q(\REGISTERS[9][20] )
         );
  DLH_X1 \REGISTERS_reg[9][19]  ( .G(n4908), .D(n5021), .Q(\REGISTERS[9][19] )
         );
  DLH_X1 \REGISTERS_reg[9][18]  ( .G(n4908), .D(n5017), .Q(\REGISTERS[9][18] )
         );
  DLH_X1 \REGISTERS_reg[9][17]  ( .G(n4908), .D(n5013), .Q(\REGISTERS[9][17] )
         );
  DLH_X1 \REGISTERS_reg[9][16]  ( .G(n4908), .D(n5008), .Q(\REGISTERS[9][16] )
         );
  DLH_X1 \REGISTERS_reg[9][15]  ( .G(n4908), .D(n5004), .Q(\REGISTERS[9][15] )
         );
  DLH_X1 \REGISTERS_reg[9][14]  ( .G(n4908), .D(n5001), .Q(\REGISTERS[9][14] )
         );
  DLH_X1 \REGISTERS_reg[9][13]  ( .G(n4908), .D(n4997), .Q(\REGISTERS[9][13] )
         );
  DLH_X1 \REGISTERS_reg[9][12]  ( .G(n4908), .D(n4993), .Q(\REGISTERS[9][12] )
         );
  DLH_X1 \REGISTERS_reg[9][11]  ( .G(n4908), .D(n4989), .Q(\REGISTERS[9][11] )
         );
  DLH_X1 \REGISTERS_reg[9][10]  ( .G(n4908), .D(n4984), .Q(\REGISTERS[9][10] )
         );
  DLH_X1 \REGISTERS_reg[9][9]  ( .G(n4910), .D(n4980), .Q(\REGISTERS[9][9] )
         );
  DLH_X1 \REGISTERS_reg[9][8]  ( .G(n4910), .D(n4977), .Q(\REGISTERS[9][8] )
         );
  DLH_X1 \REGISTERS_reg[9][7]  ( .G(n4910), .D(n4973), .Q(\REGISTERS[9][7] )
         );
  DLH_X1 \REGISTERS_reg[9][6]  ( .G(n4910), .D(n4969), .Q(\REGISTERS[9][6] )
         );
  DLH_X1 \REGISTERS_reg[9][5]  ( .G(n4910), .D(n4965), .Q(\REGISTERS[9][5] )
         );
  DLH_X1 \REGISTERS_reg[9][4]  ( .G(n4910), .D(n4962), .Q(\REGISTERS[9][4] )
         );
  DLH_X1 \REGISTERS_reg[9][3]  ( .G(n4910), .D(n4957), .Q(\REGISTERS[9][3] )
         );
  DLH_X1 \REGISTERS_reg[9][2]  ( .G(n4910), .D(n4953), .Q(\REGISTERS[9][2] )
         );
  DLH_X1 \REGISTERS_reg[9][1]  ( .G(n4910), .D(n4949), .Q(\REGISTERS[9][1] )
         );
  DLH_X1 \REGISTERS_reg[9][0]  ( .G(n4910), .D(n4944), .Q(\REGISTERS[9][0] )
         );
  DLH_X1 \REGISTERS_reg[10][31]  ( .G(n4907), .D(n5074), .Q(
        \REGISTERS[10][31] ) );
  DLH_X1 \REGISTERS_reg[10][30]  ( .G(n4907), .D(n5065), .Q(
        \REGISTERS[10][30] ) );
  DLH_X1 \REGISTERS_reg[10][29]  ( .G(n4905), .D(n5061), .Q(
        \REGISTERS[10][29] ) );
  DLH_X1 \REGISTERS_reg[10][28]  ( .G(n4905), .D(n5058), .Q(
        \REGISTERS[10][28] ) );
  DLH_X1 \REGISTERS_reg[10][27]  ( .G(n4905), .D(n5053), .Q(
        \REGISTERS[10][27] ) );
  DLH_X1 \REGISTERS_reg[10][26]  ( .G(n4905), .D(n5049), .Q(
        \REGISTERS[10][26] ) );
  DLH_X1 \REGISTERS_reg[10][25]  ( .G(n4905), .D(n5046), .Q(
        \REGISTERS[10][25] ) );
  DLH_X1 \REGISTERS_reg[10][24]  ( .G(n4905), .D(n5042), .Q(
        \REGISTERS[10][24] ) );
  DLH_X1 \REGISTERS_reg[10][23]  ( .G(n4905), .D(n5037), .Q(
        \REGISTERS[10][23] ) );
  DLH_X1 \REGISTERS_reg[10][22]  ( .G(n4905), .D(n5034), .Q(
        \REGISTERS[10][22] ) );
  DLH_X1 \REGISTERS_reg[10][21]  ( .G(n4905), .D(n5030), .Q(
        \REGISTERS[10][21] ) );
  DLH_X1 \REGISTERS_reg[10][20]  ( .G(n4905), .D(n5026), .Q(
        \REGISTERS[10][20] ) );
  DLH_X1 \REGISTERS_reg[10][19]  ( .G(n4904), .D(n5020), .Q(
        \REGISTERS[10][19] ) );
  DLH_X1 \REGISTERS_reg[10][18]  ( .G(n4904), .D(n5018), .Q(
        \REGISTERS[10][18] ) );
  DLH_X1 \REGISTERS_reg[10][17]  ( .G(n4904), .D(n5014), .Q(
        \REGISTERS[10][17] ) );
  DLH_X1 \REGISTERS_reg[10][16]  ( .G(n4904), .D(n5010), .Q(
        \REGISTERS[10][16] ) );
  DLH_X1 \REGISTERS_reg[10][15]  ( .G(n4904), .D(n5006), .Q(
        \REGISTERS[10][15] ) );
  DLH_X1 \REGISTERS_reg[10][14]  ( .G(n4904), .D(n5002), .Q(
        \REGISTERS[10][14] ) );
  DLH_X1 \REGISTERS_reg[10][13]  ( .G(n4904), .D(n4998), .Q(
        \REGISTERS[10][13] ) );
  DLH_X1 \REGISTERS_reg[10][12]  ( .G(n4904), .D(n4994), .Q(
        \REGISTERS[10][12] ) );
  DLH_X1 \REGISTERS_reg[10][11]  ( .G(n4904), .D(n4988), .Q(
        \REGISTERS[10][11] ) );
  DLH_X1 \REGISTERS_reg[10][10]  ( .G(n4904), .D(n4986), .Q(
        \REGISTERS[10][10] ) );
  DLH_X1 \REGISTERS_reg[10][9]  ( .G(n4906), .D(n4982), .Q(\REGISTERS[10][9] )
         );
  DLH_X1 \REGISTERS_reg[10][8]  ( .G(n4906), .D(n4978), .Q(\REGISTERS[10][8] )
         );
  DLH_X1 \REGISTERS_reg[10][7]  ( .G(n4906), .D(n4972), .Q(\REGISTERS[10][7] )
         );
  DLH_X1 \REGISTERS_reg[10][6]  ( .G(n4906), .D(n4970), .Q(\REGISTERS[10][6] )
         );
  DLH_X1 \REGISTERS_reg[10][5]  ( .G(n4906), .D(n4966), .Q(\REGISTERS[10][5] )
         );
  DLH_X1 \REGISTERS_reg[10][4]  ( .G(n4906), .D(n4962), .Q(\REGISTERS[10][4] )
         );
  DLH_X1 \REGISTERS_reg[10][3]  ( .G(n4906), .D(n4958), .Q(\REGISTERS[10][3] )
         );
  DLH_X1 \REGISTERS_reg[10][2]  ( .G(n4906), .D(n4954), .Q(\REGISTERS[10][2] )
         );
  DLH_X1 \REGISTERS_reg[10][1]  ( .G(n4906), .D(n4950), .Q(\REGISTERS[10][1] )
         );
  DLH_X1 \REGISTERS_reg[10][0]  ( .G(n4906), .D(n4946), .Q(\REGISTERS[10][0] )
         );
  DLH_X1 \REGISTERS_reg[11][31]  ( .G(n4903), .D(n5072), .Q(
        \REGISTERS[11][31] ) );
  DLH_X1 \REGISTERS_reg[11][30]  ( .G(n4903), .D(n5066), .Q(
        \REGISTERS[11][30] ) );
  DLH_X1 \REGISTERS_reg[11][29]  ( .G(n4901), .D(n5062), .Q(
        \REGISTERS[11][29] ) );
  DLH_X1 \REGISTERS_reg[11][28]  ( .G(n4901), .D(n5056), .Q(
        \REGISTERS[11][28] ) );
  DLH_X1 \REGISTERS_reg[11][27]  ( .G(n4901), .D(n5052), .Q(
        \REGISTERS[11][27] ) );
  DLH_X1 \REGISTERS_reg[11][26]  ( .G(n4901), .D(n5050), .Q(
        \REGISTERS[11][26] ) );
  DLH_X1 \REGISTERS_reg[11][25]  ( .G(n4901), .D(n5044), .Q(
        \REGISTERS[11][25] ) );
  DLH_X1 \REGISTERS_reg[11][24]  ( .G(n4901), .D(n5040), .Q(
        \REGISTERS[11][24] ) );
  DLH_X1 \REGISTERS_reg[11][23]  ( .G(n4901), .D(n5036), .Q(
        \REGISTERS[11][23] ) );
  DLH_X1 \REGISTERS_reg[11][22]  ( .G(n4901), .D(n5032), .Q(
        \REGISTERS[11][22] ) );
  DLH_X1 \REGISTERS_reg[11][21]  ( .G(n4901), .D(n5029), .Q(
        \REGISTERS[11][21] ) );
  DLH_X1 \REGISTERS_reg[11][20]  ( .G(n4901), .D(n5024), .Q(
        \REGISTERS[11][20] ) );
  DLH_X1 \REGISTERS_reg[11][19]  ( .G(n4900), .D(n5021), .Q(
        \REGISTERS[11][19] ) );
  DLH_X1 \REGISTERS_reg[11][18]  ( .G(n4900), .D(n5017), .Q(
        \REGISTERS[11][18] ) );
  DLH_X1 \REGISTERS_reg[11][17]  ( .G(n4900), .D(n5013), .Q(
        \REGISTERS[11][17] ) );
  DLH_X1 \REGISTERS_reg[11][16]  ( .G(n4900), .D(n5008), .Q(
        \REGISTERS[11][16] ) );
  DLH_X1 \REGISTERS_reg[11][15]  ( .G(n4900), .D(n5004), .Q(
        \REGISTERS[11][15] ) );
  DLH_X1 \REGISTERS_reg[11][14]  ( .G(n4900), .D(n5001), .Q(
        \REGISTERS[11][14] ) );
  DLH_X1 \REGISTERS_reg[11][13]  ( .G(n4900), .D(n4997), .Q(
        \REGISTERS[11][13] ) );
  DLH_X1 \REGISTERS_reg[11][12]  ( .G(n4900), .D(n4993), .Q(
        \REGISTERS[11][12] ) );
  DLH_X1 \REGISTERS_reg[11][11]  ( .G(n4900), .D(n4989), .Q(
        \REGISTERS[11][11] ) );
  DLH_X1 \REGISTERS_reg[11][10]  ( .G(n4900), .D(n4984), .Q(
        \REGISTERS[11][10] ) );
  DLH_X1 \REGISTERS_reg[11][9]  ( .G(n4902), .D(n4980), .Q(\REGISTERS[11][9] )
         );
  DLH_X1 \REGISTERS_reg[11][8]  ( .G(n4902), .D(n4977), .Q(\REGISTERS[11][8] )
         );
  DLH_X1 \REGISTERS_reg[11][7]  ( .G(n4902), .D(n4973), .Q(\REGISTERS[11][7] )
         );
  DLH_X1 \REGISTERS_reg[11][6]  ( .G(n4902), .D(n4969), .Q(\REGISTERS[11][6] )
         );
  DLH_X1 \REGISTERS_reg[11][5]  ( .G(n4902), .D(n4965), .Q(\REGISTERS[11][5] )
         );
  DLH_X1 \REGISTERS_reg[11][4]  ( .G(n4902), .D(n4960), .Q(\REGISTERS[11][4] )
         );
  DLH_X1 \REGISTERS_reg[11][3]  ( .G(n4902), .D(n4957), .Q(\REGISTERS[11][3] )
         );
  DLH_X1 \REGISTERS_reg[11][2]  ( .G(n4902), .D(n4953), .Q(\REGISTERS[11][2] )
         );
  DLH_X1 \REGISTERS_reg[11][1]  ( .G(n4902), .D(n4949), .Q(\REGISTERS[11][1] )
         );
  DLH_X1 \REGISTERS_reg[11][0]  ( .G(n4902), .D(n4945), .Q(\REGISTERS[11][0] )
         );
  DLH_X1 \REGISTERS_reg[12][31]  ( .G(n4899), .D(n5074), .Q(
        \REGISTERS[12][31] ) );
  DLH_X1 \REGISTERS_reg[12][30]  ( .G(n4899), .D(n5064), .Q(
        \REGISTERS[12][30] ) );
  DLH_X1 \REGISTERS_reg[12][29]  ( .G(n4897), .D(n5060), .Q(
        \REGISTERS[12][29] ) );
  DLH_X1 \REGISTERS_reg[12][28]  ( .G(n4897), .D(n5056), .Q(
        \REGISTERS[12][28] ) );
  DLH_X1 \REGISTERS_reg[12][27]  ( .G(n4897), .D(n5053), .Q(
        \REGISTERS[12][27] ) );
  DLH_X1 \REGISTERS_reg[12][26]  ( .G(n4897), .D(n5048), .Q(
        \REGISTERS[12][26] ) );
  DLH_X1 \REGISTERS_reg[12][25]  ( .G(n4897), .D(n5044), .Q(
        \REGISTERS[12][25] ) );
  DLH_X1 \REGISTERS_reg[12][24]  ( .G(n4897), .D(n5041), .Q(
        \REGISTERS[12][24] ) );
  DLH_X1 \REGISTERS_reg[12][23]  ( .G(n4897), .D(n5037), .Q(
        \REGISTERS[12][23] ) );
  DLH_X1 \REGISTERS_reg[12][22]  ( .G(n4897), .D(n5032), .Q(
        \REGISTERS[12][22] ) );
  DLH_X1 \REGISTERS_reg[12][21]  ( .G(n4897), .D(n5028), .Q(
        \REGISTERS[12][21] ) );
  DLH_X1 \REGISTERS_reg[12][20]  ( .G(n4897), .D(n5024), .Q(
        \REGISTERS[12][20] ) );
  DLH_X1 \REGISTERS_reg[12][19]  ( .G(n4896), .D(n5022), .Q(
        \REGISTERS[12][19] ) );
  DLH_X1 \REGISTERS_reg[12][18]  ( .G(n4896), .D(n5016), .Q(
        \REGISTERS[12][18] ) );
  DLH_X1 \REGISTERS_reg[12][17]  ( .G(n4896), .D(n5012), .Q(
        \REGISTERS[12][17] ) );
  DLH_X1 \REGISTERS_reg[12][16]  ( .G(n4896), .D(n5008), .Q(
        \REGISTERS[12][16] ) );
  DLH_X1 \REGISTERS_reg[12][15]  ( .G(n4896), .D(n5005), .Q(
        \REGISTERS[12][15] ) );
  DLH_X1 \REGISTERS_reg[12][14]  ( .G(n4896), .D(n5000), .Q(
        \REGISTERS[12][14] ) );
  DLH_X1 \REGISTERS_reg[12][13]  ( .G(n4896), .D(n4996), .Q(
        \REGISTERS[12][13] ) );
  DLH_X1 \REGISTERS_reg[12][12]  ( .G(n4896), .D(n4992), .Q(
        \REGISTERS[12][12] ) );
  DLH_X1 \REGISTERS_reg[12][11]  ( .G(n4896), .D(n4989), .Q(
        \REGISTERS[12][11] ) );
  DLH_X1 \REGISTERS_reg[12][10]  ( .G(n4896), .D(n4984), .Q(
        \REGISTERS[12][10] ) );
  DLH_X1 \REGISTERS_reg[12][9]  ( .G(n4898), .D(n4980), .Q(\REGISTERS[12][9] )
         );
  DLH_X1 \REGISTERS_reg[12][8]  ( .G(n4898), .D(n4976), .Q(\REGISTERS[12][8] )
         );
  DLH_X1 \REGISTERS_reg[12][7]  ( .G(n4898), .D(n4972), .Q(\REGISTERS[12][7] )
         );
  DLH_X1 \REGISTERS_reg[12][6]  ( .G(n4898), .D(n4968), .Q(\REGISTERS[12][6] )
         );
  DLH_X1 \REGISTERS_reg[12][5]  ( .G(n4898), .D(n4964), .Q(\REGISTERS[12][5] )
         );
  DLH_X1 \REGISTERS_reg[12][4]  ( .G(n4898), .D(n4962), .Q(\REGISTERS[12][4] )
         );
  DLH_X1 \REGISTERS_reg[12][3]  ( .G(n4898), .D(n4956), .Q(\REGISTERS[12][3] )
         );
  DLH_X1 \REGISTERS_reg[12][2]  ( .G(n4898), .D(n4952), .Q(\REGISTERS[12][2] )
         );
  DLH_X1 \REGISTERS_reg[12][1]  ( .G(n4898), .D(n4948), .Q(\REGISTERS[12][1] )
         );
  DLH_X1 \REGISTERS_reg[12][0]  ( .G(n4898), .D(n4944), .Q(\REGISTERS[12][0] )
         );
  DLH_X1 \REGISTERS_reg[13][31]  ( .G(n4895), .D(n5074), .Q(
        \REGISTERS[13][31] ) );
  DLH_X1 \REGISTERS_reg[13][30]  ( .G(n4895), .D(n5066), .Q(
        \REGISTERS[13][30] ) );
  DLH_X1 \REGISTERS_reg[13][29]  ( .G(n4893), .D(n5062), .Q(
        \REGISTERS[13][29] ) );
  DLH_X1 \REGISTERS_reg[13][28]  ( .G(n4893), .D(n5057), .Q(
        \REGISTERS[13][28] ) );
  DLH_X1 \REGISTERS_reg[13][27]  ( .G(n4893), .D(n5053), .Q(
        \REGISTERS[13][27] ) );
  DLH_X1 \REGISTERS_reg[13][26]  ( .G(n4893), .D(n5050), .Q(
        \REGISTERS[13][26] ) );
  DLH_X1 \REGISTERS_reg[13][25]  ( .G(n4893), .D(n5045), .Q(
        \REGISTERS[13][25] ) );
  DLH_X1 \REGISTERS_reg[13][24]  ( .G(n4893), .D(n5040), .Q(
        \REGISTERS[13][24] ) );
  DLH_X1 \REGISTERS_reg[13][23]  ( .G(n4893), .D(n5037), .Q(
        \REGISTERS[13][23] ) );
  DLH_X1 \REGISTERS_reg[13][22]  ( .G(n4893), .D(n5033), .Q(
        \REGISTERS[13][22] ) );
  DLH_X1 \REGISTERS_reg[13][21]  ( .G(n4893), .D(n5029), .Q(
        \REGISTERS[13][21] ) );
  DLH_X1 \REGISTERS_reg[13][20]  ( .G(n4893), .D(n5025), .Q(
        \REGISTERS[13][20] ) );
  DLH_X1 \REGISTERS_reg[13][19]  ( .G(n4892), .D(n5021), .Q(
        \REGISTERS[13][19] ) );
  DLH_X1 \REGISTERS_reg[13][18]  ( .G(n4892), .D(n5017), .Q(
        \REGISTERS[13][18] ) );
  DLH_X1 \REGISTERS_reg[13][17]  ( .G(n4892), .D(n5013), .Q(
        \REGISTERS[13][17] ) );
  DLH_X1 \REGISTERS_reg[13][16]  ( .G(n4892), .D(n5008), .Q(
        \REGISTERS[13][16] ) );
  DLH_X1 \REGISTERS_reg[13][15]  ( .G(n4892), .D(n5005), .Q(
        \REGISTERS[13][15] ) );
  DLH_X1 \REGISTERS_reg[13][14]  ( .G(n4892), .D(n5001), .Q(
        \REGISTERS[13][14] ) );
  DLH_X1 \REGISTERS_reg[13][13]  ( .G(n4892), .D(n4997), .Q(
        \REGISTERS[13][13] ) );
  DLH_X1 \REGISTERS_reg[13][12]  ( .G(n4892), .D(n4993), .Q(
        \REGISTERS[13][12] ) );
  DLH_X1 \REGISTERS_reg[13][11]  ( .G(n4892), .D(n4989), .Q(
        \REGISTERS[13][11] ) );
  DLH_X1 \REGISTERS_reg[13][10]  ( .G(n4892), .D(n4984), .Q(
        \REGISTERS[13][10] ) );
  DLH_X1 \REGISTERS_reg[13][9]  ( .G(n4894), .D(n4980), .Q(\REGISTERS[13][9] )
         );
  DLH_X1 \REGISTERS_reg[13][8]  ( .G(n4894), .D(n4977), .Q(\REGISTERS[13][8] )
         );
  DLH_X1 \REGISTERS_reg[13][7]  ( .G(n4894), .D(n4973), .Q(\REGISTERS[13][7] )
         );
  DLH_X1 \REGISTERS_reg[13][6]  ( .G(n4894), .D(n4969), .Q(\REGISTERS[13][6] )
         );
  DLH_X1 \REGISTERS_reg[13][5]  ( .G(n4894), .D(n4965), .Q(\REGISTERS[13][5] )
         );
  DLH_X1 \REGISTERS_reg[13][4]  ( .G(n4894), .D(n4962), .Q(\REGISTERS[13][4] )
         );
  DLH_X1 \REGISTERS_reg[13][3]  ( .G(n4894), .D(n4957), .Q(\REGISTERS[13][3] )
         );
  DLH_X1 \REGISTERS_reg[13][2]  ( .G(n4894), .D(n4953), .Q(\REGISTERS[13][2] )
         );
  DLH_X1 \REGISTERS_reg[13][1]  ( .G(n4894), .D(n4949), .Q(\REGISTERS[13][1] )
         );
  DLH_X1 \REGISTERS_reg[13][0]  ( .G(n4894), .D(n4945), .Q(\REGISTERS[13][0] )
         );
  DLH_X1 \REGISTERS_reg[14][31]  ( .G(n4891), .D(n5072), .Q(
        \REGISTERS[14][31] ) );
  DLH_X1 \REGISTERS_reg[14][30]  ( .G(n4891), .D(n5064), .Q(
        \REGISTERS[14][30] ) );
  DLH_X1 \REGISTERS_reg[14][29]  ( .G(n4889), .D(n5060), .Q(
        \REGISTERS[14][29] ) );
  DLH_X1 \REGISTERS_reg[14][28]  ( .G(n4889), .D(n5056), .Q(
        \REGISTERS[14][28] ) );
  DLH_X1 \REGISTERS_reg[14][27]  ( .G(n4889), .D(n5053), .Q(
        \REGISTERS[14][27] ) );
  DLH_X1 \REGISTERS_reg[14][26]  ( .G(n4889), .D(n5048), .Q(
        \REGISTERS[14][26] ) );
  DLH_X1 \REGISTERS_reg[14][25]  ( .G(n4889), .D(n5044), .Q(
        \REGISTERS[14][25] ) );
  DLH_X1 \REGISTERS_reg[14][24]  ( .G(n4889), .D(n5040), .Q(
        \REGISTERS[14][24] ) );
  DLH_X1 \REGISTERS_reg[14][23]  ( .G(n4889), .D(n5037), .Q(
        \REGISTERS[14][23] ) );
  DLH_X1 \REGISTERS_reg[14][22]  ( .G(n4889), .D(n5032), .Q(
        \REGISTERS[14][22] ) );
  DLH_X1 \REGISTERS_reg[14][21]  ( .G(n4889), .D(n5028), .Q(
        \REGISTERS[14][21] ) );
  DLH_X1 \REGISTERS_reg[14][20]  ( .G(n4889), .D(n5024), .Q(
        \REGISTERS[14][20] ) );
  DLH_X1 \REGISTERS_reg[14][19]  ( .G(n4888), .D(n5022), .Q(
        \REGISTERS[14][19] ) );
  DLH_X1 \REGISTERS_reg[14][18]  ( .G(n4888), .D(n5016), .Q(
        \REGISTERS[14][18] ) );
  DLH_X1 \REGISTERS_reg[14][17]  ( .G(n4888), .D(n5012), .Q(
        \REGISTERS[14][17] ) );
  DLH_X1 \REGISTERS_reg[14][16]  ( .G(n4888), .D(n5008), .Q(
        \REGISTERS[14][16] ) );
  DLH_X1 \REGISTERS_reg[14][15]  ( .G(n4888), .D(n5005), .Q(
        \REGISTERS[14][15] ) );
  DLH_X1 \REGISTERS_reg[14][14]  ( .G(n4888), .D(n5000), .Q(
        \REGISTERS[14][14] ) );
  DLH_X1 \REGISTERS_reg[14][13]  ( .G(n4888), .D(n4996), .Q(
        \REGISTERS[14][13] ) );
  DLH_X1 \REGISTERS_reg[14][12]  ( .G(n4888), .D(n4992), .Q(
        \REGISTERS[14][12] ) );
  DLH_X1 \REGISTERS_reg[14][11]  ( .G(n4888), .D(n4989), .Q(
        \REGISTERS[14][11] ) );
  DLH_X1 \REGISTERS_reg[14][10]  ( .G(n4888), .D(n4984), .Q(
        \REGISTERS[14][10] ) );
  DLH_X1 \REGISTERS_reg[14][9]  ( .G(n4890), .D(n4980), .Q(\REGISTERS[14][9] )
         );
  DLH_X1 \REGISTERS_reg[14][8]  ( .G(n4890), .D(n4976), .Q(\REGISTERS[14][8] )
         );
  DLH_X1 \REGISTERS_reg[14][7]  ( .G(n4890), .D(n4972), .Q(\REGISTERS[14][7] )
         );
  DLH_X1 \REGISTERS_reg[14][6]  ( .G(n4890), .D(n4968), .Q(\REGISTERS[14][6] )
         );
  DLH_X1 \REGISTERS_reg[14][5]  ( .G(n4890), .D(n4964), .Q(\REGISTERS[14][5] )
         );
  DLH_X1 \REGISTERS_reg[14][4]  ( .G(n4890), .D(n4960), .Q(\REGISTERS[14][4] )
         );
  DLH_X1 \REGISTERS_reg[14][3]  ( .G(n4890), .D(n4956), .Q(\REGISTERS[14][3] )
         );
  DLH_X1 \REGISTERS_reg[14][2]  ( .G(n4890), .D(n4952), .Q(\REGISTERS[14][2] )
         );
  DLH_X1 \REGISTERS_reg[14][1]  ( .G(n4890), .D(n4948), .Q(\REGISTERS[14][1] )
         );
  DLH_X1 \REGISTERS_reg[14][0]  ( .G(n4890), .D(n4944), .Q(\REGISTERS[14][0] )
         );
  DLH_X1 \REGISTERS_reg[15][31]  ( .G(n4887), .D(n5073), .Q(
        \REGISTERS[15][31] ) );
  DLH_X1 \REGISTERS_reg[15][30]  ( .G(n4887), .D(n5065), .Q(
        \REGISTERS[15][30] ) );
  DLH_X1 \REGISTERS_reg[15][29]  ( .G(n4885), .D(n5061), .Q(
        \REGISTERS[15][29] ) );
  DLH_X1 \REGISTERS_reg[15][28]  ( .G(n4885), .D(n5058), .Q(
        \REGISTERS[15][28] ) );
  DLH_X1 \REGISTERS_reg[15][27]  ( .G(n4885), .D(n5052), .Q(
        \REGISTERS[15][27] ) );
  DLH_X1 \REGISTERS_reg[15][26]  ( .G(n4885), .D(n5049), .Q(
        \REGISTERS[15][26] ) );
  DLH_X1 \REGISTERS_reg[15][25]  ( .G(n4885), .D(n5046), .Q(
        \REGISTERS[15][25] ) );
  DLH_X1 \REGISTERS_reg[15][24]  ( .G(n4885), .D(n5042), .Q(
        \REGISTERS[15][24] ) );
  DLH_X1 \REGISTERS_reg[15][23]  ( .G(n4885), .D(n5036), .Q(
        \REGISTERS[15][23] ) );
  DLH_X1 \REGISTERS_reg[15][22]  ( .G(n4885), .D(n5034), .Q(
        \REGISTERS[15][22] ) );
  DLH_X1 \REGISTERS_reg[15][21]  ( .G(n4885), .D(n5030), .Q(
        \REGISTERS[15][21] ) );
  DLH_X1 \REGISTERS_reg[15][20]  ( .G(n4885), .D(n5026), .Q(
        \REGISTERS[15][20] ) );
  DLH_X1 \REGISTERS_reg[15][19]  ( .G(n4884), .D(n5021), .Q(
        \REGISTERS[15][19] ) );
  DLH_X1 \REGISTERS_reg[15][18]  ( .G(n4884), .D(n5018), .Q(
        \REGISTERS[15][18] ) );
  DLH_X1 \REGISTERS_reg[15][17]  ( .G(n4884), .D(n5014), .Q(
        \REGISTERS[15][17] ) );
  DLH_X1 \REGISTERS_reg[15][16]  ( .G(n4884), .D(n5010), .Q(
        \REGISTERS[15][16] ) );
  DLH_X1 \REGISTERS_reg[15][15]  ( .G(n4884), .D(n5006), .Q(
        \REGISTERS[15][15] ) );
  DLH_X1 \REGISTERS_reg[15][14]  ( .G(n4884), .D(n5002), .Q(
        \REGISTERS[15][14] ) );
  DLH_X1 \REGISTERS_reg[15][13]  ( .G(n4884), .D(n4998), .Q(
        \REGISTERS[15][13] ) );
  DLH_X1 \REGISTERS_reg[15][12]  ( .G(n4884), .D(n4994), .Q(
        \REGISTERS[15][12] ) );
  DLH_X1 \REGISTERS_reg[15][11]  ( .G(n4884), .D(n4988), .Q(
        \REGISTERS[15][11] ) );
  DLH_X1 \REGISTERS_reg[15][10]  ( .G(n4884), .D(n4986), .Q(
        \REGISTERS[15][10] ) );
  DLH_X1 \REGISTERS_reg[15][9]  ( .G(n4886), .D(n4982), .Q(\REGISTERS[15][9] )
         );
  DLH_X1 \REGISTERS_reg[15][8]  ( .G(n4886), .D(n4978), .Q(\REGISTERS[15][8] )
         );
  DLH_X1 \REGISTERS_reg[15][7]  ( .G(n4886), .D(n4973), .Q(\REGISTERS[15][7] )
         );
  DLH_X1 \REGISTERS_reg[15][6]  ( .G(n4886), .D(n4970), .Q(\REGISTERS[15][6] )
         );
  DLH_X1 \REGISTERS_reg[15][5]  ( .G(n4886), .D(n4966), .Q(\REGISTERS[15][5] )
         );
  DLH_X1 \REGISTERS_reg[15][4]  ( .G(n4886), .D(n4962), .Q(\REGISTERS[15][4] )
         );
  DLH_X1 \REGISTERS_reg[15][3]  ( .G(n4886), .D(n4958), .Q(\REGISTERS[15][3] )
         );
  DLH_X1 \REGISTERS_reg[15][2]  ( .G(n4886), .D(n4954), .Q(\REGISTERS[15][2] )
         );
  DLH_X1 \REGISTERS_reg[15][1]  ( .G(n4886), .D(n4950), .Q(\REGISTERS[15][1] )
         );
  DLH_X1 \REGISTERS_reg[15][0]  ( .G(n4886), .D(n4946), .Q(\REGISTERS[15][0] )
         );
  DLH_X1 \REGISTERS_reg[16][31]  ( .G(n4883), .D(n5072), .Q(
        \REGISTERS[16][31] ) );
  DLH_X1 \REGISTERS_reg[16][30]  ( .G(n4883), .D(n5067), .Q(
        \REGISTERS[16][30] ) );
  DLH_X1 \REGISTERS_reg[16][29]  ( .G(n4881), .D(n5063), .Q(
        \REGISTERS[16][29] ) );
  DLH_X1 \REGISTERS_reg[16][28]  ( .G(n4881), .D(n5059), .Q(
        \REGISTERS[16][28] ) );
  DLH_X1 \REGISTERS_reg[16][27]  ( .G(n4881), .D(n5054), .Q(
        \REGISTERS[16][27] ) );
  DLH_X1 \REGISTERS_reg[16][26]  ( .G(n4881), .D(n5051), .Q(
        \REGISTERS[16][26] ) );
  DLH_X1 \REGISTERS_reg[16][25]  ( .G(n4881), .D(n5047), .Q(
        \REGISTERS[16][25] ) );
  DLH_X1 \REGISTERS_reg[16][24]  ( .G(n4881), .D(n5040), .Q(
        \REGISTERS[16][24] ) );
  DLH_X1 \REGISTERS_reg[16][23]  ( .G(n4881), .D(n5038), .Q(
        \REGISTERS[16][23] ) );
  DLH_X1 \REGISTERS_reg[16][22]  ( .G(n4881), .D(n5035), .Q(
        \REGISTERS[16][22] ) );
  DLH_X1 \REGISTERS_reg[16][21]  ( .G(n4881), .D(n5030), .Q(
        \REGISTERS[16][21] ) );
  DLH_X1 \REGISTERS_reg[16][20]  ( .G(n4881), .D(n5027), .Q(
        \REGISTERS[16][20] ) );
  DLH_X1 \REGISTERS_reg[16][19]  ( .G(n4880), .D(n5022), .Q(
        \REGISTERS[16][19] ) );
  DLH_X1 \REGISTERS_reg[16][18]  ( .G(n4880), .D(n5018), .Q(
        \REGISTERS[16][18] ) );
  DLH_X1 \REGISTERS_reg[16][17]  ( .G(n4880), .D(n5014), .Q(
        \REGISTERS[16][17] ) );
  DLH_X1 \REGISTERS_reg[16][16]  ( .G(n4880), .D(n5010), .Q(
        \REGISTERS[16][16] ) );
  DLH_X1 \REGISTERS_reg[16][15]  ( .G(n4880), .D(n5007), .Q(
        \REGISTERS[16][15] ) );
  DLH_X1 \REGISTERS_reg[16][14]  ( .G(n4880), .D(n5002), .Q(
        \REGISTERS[16][14] ) );
  DLH_X1 \REGISTERS_reg[16][13]  ( .G(n4880), .D(n4998), .Q(
        \REGISTERS[16][13] ) );
  DLH_X1 \REGISTERS_reg[16][12]  ( .G(n4880), .D(n4994), .Q(
        \REGISTERS[16][12] ) );
  DLH_X1 \REGISTERS_reg[16][11]  ( .G(n4880), .D(n4990), .Q(
        \REGISTERS[16][11] ) );
  DLH_X1 \REGISTERS_reg[16][10]  ( .G(n4880), .D(n4986), .Q(
        \REGISTERS[16][10] ) );
  DLH_X1 \REGISTERS_reg[16][9]  ( .G(n4882), .D(n4982), .Q(\REGISTERS[16][9] )
         );
  DLH_X1 \REGISTERS_reg[16][8]  ( .G(n4882), .D(n4978), .Q(\REGISTERS[16][8] )
         );
  DLH_X1 \REGISTERS_reg[16][7]  ( .G(n4882), .D(n4974), .Q(\REGISTERS[16][7] )
         );
  DLH_X1 \REGISTERS_reg[16][6]  ( .G(n4882), .D(n4970), .Q(\REGISTERS[16][6] )
         );
  DLH_X1 \REGISTERS_reg[16][5]  ( .G(n4882), .D(n4966), .Q(\REGISTERS[16][5] )
         );
  DLH_X1 \REGISTERS_reg[16][4]  ( .G(n4882), .D(n4960), .Q(\REGISTERS[16][4] )
         );
  DLH_X1 \REGISTERS_reg[16][3]  ( .G(n4882), .D(n4958), .Q(\REGISTERS[16][3] )
         );
  DLH_X1 \REGISTERS_reg[16][2]  ( .G(n4882), .D(n4954), .Q(\REGISTERS[16][2] )
         );
  DLH_X1 \REGISTERS_reg[16][1]  ( .G(n4882), .D(n4950), .Q(\REGISTERS[16][1] )
         );
  DLH_X1 \REGISTERS_reg[16][0]  ( .G(n4882), .D(n4946), .Q(\REGISTERS[16][0] )
         );
  DLH_X1 \REGISTERS_reg[17][31]  ( .G(n4879), .D(n5073), .Q(
        \REGISTERS[17][31] ) );
  DLH_X1 \REGISTERS_reg[17][30]  ( .G(n4879), .D(n5064), .Q(
        \REGISTERS[17][30] ) );
  DLH_X1 \REGISTERS_reg[17][29]  ( .G(n4877), .D(n5060), .Q(
        \REGISTERS[17][29] ) );
  DLH_X1 \REGISTERS_reg[17][28]  ( .G(n4877), .D(n5056), .Q(
        \REGISTERS[17][28] ) );
  DLH_X1 \REGISTERS_reg[17][27]  ( .G(n4877), .D(n5052), .Q(
        \REGISTERS[17][27] ) );
  DLH_X1 \REGISTERS_reg[17][26]  ( .G(n4877), .D(n5048), .Q(
        \REGISTERS[17][26] ) );
  DLH_X1 \REGISTERS_reg[17][25]  ( .G(n4877), .D(n5044), .Q(
        \REGISTERS[17][25] ) );
  DLH_X1 \REGISTERS_reg[17][24]  ( .G(n4877), .D(n5041), .Q(
        \REGISTERS[17][24] ) );
  DLH_X1 \REGISTERS_reg[17][23]  ( .G(n4877), .D(n5036), .Q(
        \REGISTERS[17][23] ) );
  DLH_X1 \REGISTERS_reg[17][22]  ( .G(n4877), .D(n5032), .Q(
        \REGISTERS[17][22] ) );
  DLH_X1 \REGISTERS_reg[17][21]  ( .G(n4877), .D(n5029), .Q(
        \REGISTERS[17][21] ) );
  DLH_X1 \REGISTERS_reg[17][20]  ( .G(n4877), .D(n5024), .Q(
        \REGISTERS[17][20] ) );
  DLH_X1 \REGISTERS_reg[17][19]  ( .G(n4876), .D(n5023), .Q(
        \REGISTERS[17][19] ) );
  DLH_X1 \REGISTERS_reg[17][18]  ( .G(n4876), .D(n5017), .Q(
        \REGISTERS[17][18] ) );
  DLH_X1 \REGISTERS_reg[17][17]  ( .G(n4876), .D(n5015), .Q(
        \REGISTERS[17][17] ) );
  DLH_X1 \REGISTERS_reg[17][16]  ( .G(n4876), .D(n5009), .Q(
        \REGISTERS[17][16] ) );
  DLH_X1 \REGISTERS_reg[17][15]  ( .G(n4876), .D(n5004), .Q(
        \REGISTERS[17][15] ) );
  DLH_X1 \REGISTERS_reg[17][14]  ( .G(n4876), .D(n5001), .Q(
        \REGISTERS[17][14] ) );
  DLH_X1 \REGISTERS_reg[17][13]  ( .G(n4876), .D(n4996), .Q(
        \REGISTERS[17][13] ) );
  DLH_X1 \REGISTERS_reg[17][12]  ( .G(n4876), .D(n4995), .Q(
        \REGISTERS[17][12] ) );
  DLH_X1 \REGISTERS_reg[17][11]  ( .G(n4876), .D(n4991), .Q(
        \REGISTERS[17][11] ) );
  DLH_X1 \REGISTERS_reg[17][10]  ( .G(n4876), .D(n4985), .Q(
        \REGISTERS[17][10] ) );
  DLH_X1 \REGISTERS_reg[17][9]  ( .G(n4878), .D(n4981), .Q(\REGISTERS[17][9] )
         );
  DLH_X1 \REGISTERS_reg[17][8]  ( .G(n4878), .D(n4979), .Q(\REGISTERS[17][8] )
         );
  DLH_X1 \REGISTERS_reg[17][7]  ( .G(n4878), .D(n4973), .Q(\REGISTERS[17][7] )
         );
  DLH_X1 \REGISTERS_reg[17][6]  ( .G(n4878), .D(n4971), .Q(\REGISTERS[17][6] )
         );
  DLH_X1 \REGISTERS_reg[17][5]  ( .G(n4878), .D(n4967), .Q(\REGISTERS[17][5] )
         );
  DLH_X1 \REGISTERS_reg[17][4]  ( .G(n4878), .D(n4961), .Q(\REGISTERS[17][4] )
         );
  DLH_X1 \REGISTERS_reg[17][3]  ( .G(n4878), .D(n4957), .Q(\REGISTERS[17][3] )
         );
  DLH_X1 \REGISTERS_reg[17][2]  ( .G(n4878), .D(n4953), .Q(\REGISTERS[17][2] )
         );
  DLH_X1 \REGISTERS_reg[17][1]  ( .G(n4878), .D(n4948), .Q(\REGISTERS[17][1] )
         );
  DLH_X1 \REGISTERS_reg[17][0]  ( .G(n4878), .D(n4947), .Q(\REGISTERS[17][0] )
         );
  DLH_X1 \REGISTERS_reg[18][31]  ( .G(n4875), .D(n5074), .Q(
        \REGISTERS[18][31] ) );
  DLH_X1 \REGISTERS_reg[18][30]  ( .G(n4875), .D(n5067), .Q(
        \REGISTERS[18][30] ) );
  DLH_X1 \REGISTERS_reg[18][29]  ( .G(n4873), .D(n5063), .Q(
        \REGISTERS[18][29] ) );
  DLH_X1 \REGISTERS_reg[18][28]  ( .G(n4873), .D(n5059), .Q(
        \REGISTERS[18][28] ) );
  DLH_X1 \REGISTERS_reg[18][27]  ( .G(n4873), .D(n5055), .Q(
        \REGISTERS[18][27] ) );
  DLH_X1 \REGISTERS_reg[18][26]  ( .G(n4873), .D(n5051), .Q(
        \REGISTERS[18][26] ) );
  DLH_X1 \REGISTERS_reg[18][25]  ( .G(n4873), .D(n5047), .Q(
        \REGISTERS[18][25] ) );
  DLH_X1 \REGISTERS_reg[18][24]  ( .G(n4873), .D(n5043), .Q(
        \REGISTERS[18][24] ) );
  DLH_X1 \REGISTERS_reg[18][23]  ( .G(n4873), .D(n5039), .Q(
        \REGISTERS[18][23] ) );
  DLH_X1 \REGISTERS_reg[18][22]  ( .G(n4873), .D(n5035), .Q(
        \REGISTERS[18][22] ) );
  DLH_X1 \REGISTERS_reg[18][21]  ( .G(n4873), .D(n5030), .Q(
        \REGISTERS[18][21] ) );
  DLH_X1 \REGISTERS_reg[18][20]  ( .G(n4873), .D(n5027), .Q(
        \REGISTERS[18][20] ) );
  DLH_X1 \REGISTERS_reg[18][19]  ( .G(n4872), .D(n5022), .Q(
        \REGISTERS[18][19] ) );
  DLH_X1 \REGISTERS_reg[18][18]  ( .G(n4872), .D(n5018), .Q(
        \REGISTERS[18][18] ) );
  DLH_X1 \REGISTERS_reg[18][17]  ( .G(n4872), .D(n5012), .Q(
        \REGISTERS[18][17] ) );
  DLH_X1 \REGISTERS_reg[18][16]  ( .G(n4872), .D(n5010), .Q(
        \REGISTERS[18][16] ) );
  DLH_X1 \REGISTERS_reg[18][15]  ( .G(n4872), .D(n5007), .Q(
        \REGISTERS[18][15] ) );
  DLH_X1 \REGISTERS_reg[18][14]  ( .G(n4872), .D(n5002), .Q(
        \REGISTERS[18][14] ) );
  DLH_X1 \REGISTERS_reg[18][13]  ( .G(n4872), .D(n4999), .Q(
        \REGISTERS[18][13] ) );
  DLH_X1 \REGISTERS_reg[18][12]  ( .G(n4872), .D(n4992), .Q(
        \REGISTERS[18][12] ) );
  DLH_X1 \REGISTERS_reg[18][11]  ( .G(n4872), .D(n4991), .Q(
        \REGISTERS[18][11] ) );
  DLH_X1 \REGISTERS_reg[18][10]  ( .G(n4872), .D(n4986), .Q(
        \REGISTERS[18][10] ) );
  DLH_X1 \REGISTERS_reg[18][9]  ( .G(n4874), .D(n4982), .Q(\REGISTERS[18][9] )
         );
  DLH_X1 \REGISTERS_reg[18][8]  ( .G(n4874), .D(n4976), .Q(\REGISTERS[18][8] )
         );
  DLH_X1 \REGISTERS_reg[18][7]  ( .G(n4874), .D(n4974), .Q(\REGISTERS[18][7] )
         );
  DLH_X1 \REGISTERS_reg[18][6]  ( .G(n4874), .D(n4968), .Q(\REGISTERS[18][6] )
         );
  DLH_X1 \REGISTERS_reg[18][5]  ( .G(n4874), .D(n4964), .Q(\REGISTERS[18][5] )
         );
  DLH_X1 \REGISTERS_reg[18][4]  ( .G(n4874), .D(n4962), .Q(\REGISTERS[18][4] )
         );
  DLH_X1 \REGISTERS_reg[18][3]  ( .G(n4874), .D(n4958), .Q(\REGISTERS[18][3] )
         );
  DLH_X1 \REGISTERS_reg[18][2]  ( .G(n4874), .D(n4954), .Q(\REGISTERS[18][2] )
         );
  DLH_X1 \REGISTERS_reg[18][1]  ( .G(n4874), .D(n4951), .Q(\REGISTERS[18][1] )
         );
  DLH_X1 \REGISTERS_reg[18][0]  ( .G(n4874), .D(n4944), .Q(\REGISTERS[18][0] )
         );
  DLH_X1 \REGISTERS_reg[19][31]  ( .G(n4871), .D(n5073), .Q(
        \REGISTERS[19][31] ) );
  DLH_X1 \REGISTERS_reg[19][30]  ( .G(n4871), .D(n5066), .Q(
        \REGISTERS[19][30] ) );
  DLH_X1 \REGISTERS_reg[19][29]  ( .G(n4869), .D(n5062), .Q(
        \REGISTERS[19][29] ) );
  DLH_X1 \REGISTERS_reg[19][28]  ( .G(n4869), .D(n5058), .Q(
        \REGISTERS[19][28] ) );
  DLH_X1 \REGISTERS_reg[19][27]  ( .G(n4869), .D(n5054), .Q(
        \REGISTERS[19][27] ) );
  DLH_X1 \REGISTERS_reg[19][26]  ( .G(n4869), .D(n5050), .Q(
        \REGISTERS[19][26] ) );
  DLH_X1 \REGISTERS_reg[19][25]  ( .G(n4869), .D(n5046), .Q(
        \REGISTERS[19][25] ) );
  DLH_X1 \REGISTERS_reg[19][24]  ( .G(n4869), .D(n5041), .Q(
        \REGISTERS[19][24] ) );
  DLH_X1 \REGISTERS_reg[19][23]  ( .G(n4869), .D(n5038), .Q(
        \REGISTERS[19][23] ) );
  DLH_X1 \REGISTERS_reg[19][22]  ( .G(n4869), .D(n5034), .Q(
        \REGISTERS[19][22] ) );
  DLH_X1 \REGISTERS_reg[19][21]  ( .G(n4869), .D(n5029), .Q(
        \REGISTERS[19][21] ) );
  DLH_X1 \REGISTERS_reg[19][20]  ( .G(n4869), .D(n5026), .Q(
        \REGISTERS[19][20] ) );
  DLH_X1 \REGISTERS_reg[19][19]  ( .G(n4868), .D(n5021), .Q(
        \REGISTERS[19][19] ) );
  DLH_X1 \REGISTERS_reg[19][18]  ( .G(n4868), .D(n5017), .Q(
        \REGISTERS[19][18] ) );
  DLH_X1 \REGISTERS_reg[19][17]  ( .G(n4868), .D(n5013), .Q(
        \REGISTERS[19][17] ) );
  DLH_X1 \REGISTERS_reg[19][16]  ( .G(n4868), .D(n5009), .Q(
        \REGISTERS[19][16] ) );
  DLH_X1 \REGISTERS_reg[19][15]  ( .G(n4868), .D(n5004), .Q(
        \REGISTERS[19][15] ) );
  DLH_X1 \REGISTERS_reg[19][14]  ( .G(n4868), .D(n5001), .Q(
        \REGISTERS[19][14] ) );
  DLH_X1 \REGISTERS_reg[19][13]  ( .G(n4868), .D(n4998), .Q(
        \REGISTERS[19][13] ) );
  DLH_X1 \REGISTERS_reg[19][12]  ( .G(n4868), .D(n4993), .Q(
        \REGISTERS[19][12] ) );
  DLH_X1 \REGISTERS_reg[19][11]  ( .G(n4868), .D(n4990), .Q(
        \REGISTERS[19][11] ) );
  DLH_X1 \REGISTERS_reg[19][10]  ( .G(n4868), .D(n4985), .Q(
        \REGISTERS[19][10] ) );
  DLH_X1 \REGISTERS_reg[19][9]  ( .G(n4870), .D(n4981), .Q(\REGISTERS[19][9] )
         );
  DLH_X1 \REGISTERS_reg[19][8]  ( .G(n4870), .D(n4977), .Q(\REGISTERS[19][8] )
         );
  DLH_X1 \REGISTERS_reg[19][7]  ( .G(n4870), .D(n4973), .Q(\REGISTERS[19][7] )
         );
  DLH_X1 \REGISTERS_reg[19][6]  ( .G(n4870), .D(n4969), .Q(\REGISTERS[19][6] )
         );
  DLH_X1 \REGISTERS_reg[19][5]  ( .G(n4870), .D(n4965), .Q(\REGISTERS[19][5] )
         );
  DLH_X1 \REGISTERS_reg[19][4]  ( .G(n4870), .D(n4961), .Q(\REGISTERS[19][4] )
         );
  DLH_X1 \REGISTERS_reg[19][3]  ( .G(n4870), .D(n4957), .Q(\REGISTERS[19][3] )
         );
  DLH_X1 \REGISTERS_reg[19][2]  ( .G(n4870), .D(n4953), .Q(\REGISTERS[19][2] )
         );
  DLH_X1 \REGISTERS_reg[19][1]  ( .G(n4870), .D(n4950), .Q(\REGISTERS[19][1] )
         );
  DLH_X1 \REGISTERS_reg[19][0]  ( .G(n4870), .D(n4946), .Q(\REGISTERS[19][0] )
         );
  DLH_X1 \REGISTERS_reg[20][31]  ( .G(n4867), .D(n5075), .Q(
        \REGISTERS[20][31] ) );
  DLH_X1 \REGISTERS_reg[20][30]  ( .G(n4867), .D(n5064), .Q(
        \REGISTERS[20][30] ) );
  DLH_X1 \REGISTERS_reg[20][29]  ( .G(n4865), .D(n5060), .Q(
        \REGISTERS[20][29] ) );
  DLH_X1 \REGISTERS_reg[20][28]  ( .G(n4865), .D(n5056), .Q(
        \REGISTERS[20][28] ) );
  DLH_X1 \REGISTERS_reg[20][27]  ( .G(n4865), .D(n5052), .Q(
        \REGISTERS[20][27] ) );
  DLH_X1 \REGISTERS_reg[20][26]  ( .G(n4865), .D(n5048), .Q(
        \REGISTERS[20][26] ) );
  DLH_X1 \REGISTERS_reg[20][25]  ( .G(n4865), .D(n5044), .Q(
        \REGISTERS[20][25] ) );
  DLH_X1 \REGISTERS_reg[20][24]  ( .G(n4865), .D(n5042), .Q(
        \REGISTERS[20][24] ) );
  DLH_X1 \REGISTERS_reg[20][23]  ( .G(n4865), .D(n5036), .Q(
        \REGISTERS[20][23] ) );
  DLH_X1 \REGISTERS_reg[20][22]  ( .G(n4865), .D(n5032), .Q(
        \REGISTERS[20][22] ) );
  DLH_X1 \REGISTERS_reg[20][21]  ( .G(n4865), .D(n5028), .Q(
        \REGISTERS[20][21] ) );
  DLH_X1 \REGISTERS_reg[20][20]  ( .G(n4865), .D(n5024), .Q(
        \REGISTERS[20][20] ) );
  DLH_X1 \REGISTERS_reg[20][19]  ( .G(n4864), .D(n5020), .Q(
        \REGISTERS[20][19] ) );
  DLH_X1 \REGISTERS_reg[20][18]  ( .G(n4864), .D(n5016), .Q(
        \REGISTERS[20][18] ) );
  DLH_X1 \REGISTERS_reg[20][17]  ( .G(n4864), .D(n5012), .Q(
        \REGISTERS[20][17] ) );
  DLH_X1 \REGISTERS_reg[20][16]  ( .G(n4864), .D(n5009), .Q(
        \REGISTERS[20][16] ) );
  DLH_X1 \REGISTERS_reg[20][15]  ( .G(n4864), .D(n5004), .Q(
        \REGISTERS[20][15] ) );
  DLH_X1 \REGISTERS_reg[20][14]  ( .G(n4864), .D(n5000), .Q(
        \REGISTERS[20][14] ) );
  DLH_X1 \REGISTERS_reg[20][13]  ( .G(n4864), .D(n4996), .Q(
        \REGISTERS[20][13] ) );
  DLH_X1 \REGISTERS_reg[20][12]  ( .G(n4864), .D(n4992), .Q(
        \REGISTERS[20][12] ) );
  DLH_X1 \REGISTERS_reg[20][11]  ( .G(n4864), .D(n4988), .Q(
        \REGISTERS[20][11] ) );
  DLH_X1 \REGISTERS_reg[20][10]  ( .G(n4864), .D(n4985), .Q(
        \REGISTERS[20][10] ) );
  DLH_X1 \REGISTERS_reg[20][9]  ( .G(n4866), .D(n4981), .Q(\REGISTERS[20][9] )
         );
  DLH_X1 \REGISTERS_reg[20][8]  ( .G(n4866), .D(n4976), .Q(\REGISTERS[20][8] )
         );
  DLH_X1 \REGISTERS_reg[20][7]  ( .G(n4866), .D(n4972), .Q(\REGISTERS[20][7] )
         );
  DLH_X1 \REGISTERS_reg[20][6]  ( .G(n4866), .D(n4968), .Q(\REGISTERS[20][6] )
         );
  DLH_X1 \REGISTERS_reg[20][5]  ( .G(n4866), .D(n4964), .Q(\REGISTERS[20][5] )
         );
  DLH_X1 \REGISTERS_reg[20][4]  ( .G(n4866), .D(n4962), .Q(\REGISTERS[20][4] )
         );
  DLH_X1 \REGISTERS_reg[20][3]  ( .G(n4866), .D(n4956), .Q(\REGISTERS[20][3] )
         );
  DLH_X1 \REGISTERS_reg[20][2]  ( .G(n4866), .D(n4952), .Q(\REGISTERS[20][2] )
         );
  DLH_X1 \REGISTERS_reg[20][1]  ( .G(n4866), .D(n4948), .Q(\REGISTERS[20][1] )
         );
  DLH_X1 \REGISTERS_reg[20][0]  ( .G(n4866), .D(n4944), .Q(\REGISTERS[20][0] )
         );
  DLH_X1 \REGISTERS_reg[21][31]  ( .G(n4863), .D(n5075), .Q(
        \REGISTERS[21][31] ) );
  DLH_X1 \REGISTERS_reg[21][30]  ( .G(n4863), .D(n5066), .Q(
        \REGISTERS[21][30] ) );
  DLH_X1 \REGISTERS_reg[21][29]  ( .G(n4861), .D(n5062), .Q(
        \REGISTERS[21][29] ) );
  DLH_X1 \REGISTERS_reg[21][28]  ( .G(n4861), .D(n5058), .Q(
        \REGISTERS[21][28] ) );
  DLH_X1 \REGISTERS_reg[21][27]  ( .G(n4861), .D(n5054), .Q(
        \REGISTERS[21][27] ) );
  DLH_X1 \REGISTERS_reg[21][26]  ( .G(n4861), .D(n5050), .Q(
        \REGISTERS[21][26] ) );
  DLH_X1 \REGISTERS_reg[21][25]  ( .G(n4861), .D(n5046), .Q(
        \REGISTERS[21][25] ) );
  DLH_X1 \REGISTERS_reg[21][24]  ( .G(n4861), .D(n5042), .Q(
        \REGISTERS[21][24] ) );
  DLH_X1 \REGISTERS_reg[21][23]  ( .G(n4861), .D(n5038), .Q(
        \REGISTERS[21][23] ) );
  DLH_X1 \REGISTERS_reg[21][22]  ( .G(n4861), .D(n5034), .Q(
        \REGISTERS[21][22] ) );
  DLH_X1 \REGISTERS_reg[21][21]  ( .G(n4861), .D(n5028), .Q(
        \REGISTERS[21][21] ) );
  DLH_X1 \REGISTERS_reg[21][20]  ( .G(n4861), .D(n5026), .Q(
        \REGISTERS[21][20] ) );
  DLH_X1 \REGISTERS_reg[21][19]  ( .G(n4860), .D(n5021), .Q(
        \REGISTERS[21][19] ) );
  DLH_X1 \REGISTERS_reg[21][18]  ( .G(n4860), .D(n5016), .Q(
        \REGISTERS[21][18] ) );
  DLH_X1 \REGISTERS_reg[21][17]  ( .G(n4860), .D(n5013), .Q(
        \REGISTERS[21][17] ) );
  DLH_X1 \REGISTERS_reg[21][16]  ( .G(n4860), .D(n5009), .Q(
        \REGISTERS[21][16] ) );
  DLH_X1 \REGISTERS_reg[21][15]  ( .G(n4860), .D(n5004), .Q(
        \REGISTERS[21][15] ) );
  DLH_X1 \REGISTERS_reg[21][14]  ( .G(n4860), .D(n5000), .Q(
        \REGISTERS[21][14] ) );
  DLH_X1 \REGISTERS_reg[21][13]  ( .G(n4860), .D(n4996), .Q(
        \REGISTERS[21][13] ) );
  DLH_X1 \REGISTERS_reg[21][12]  ( .G(n4860), .D(n4993), .Q(
        \REGISTERS[21][12] ) );
  DLH_X1 \REGISTERS_reg[21][11]  ( .G(n4860), .D(n4990), .Q(
        \REGISTERS[21][11] ) );
  DLH_X1 \REGISTERS_reg[21][10]  ( .G(n4860), .D(n4985), .Q(
        \REGISTERS[21][10] ) );
  DLH_X1 \REGISTERS_reg[21][9]  ( .G(n4862), .D(n4981), .Q(\REGISTERS[21][9] )
         );
  DLH_X1 \REGISTERS_reg[21][8]  ( .G(n4862), .D(n4977), .Q(\REGISTERS[21][8] )
         );
  DLH_X1 \REGISTERS_reg[21][7]  ( .G(n4862), .D(n4975), .Q(\REGISTERS[21][7] )
         );
  DLH_X1 \REGISTERS_reg[21][6]  ( .G(n4862), .D(n4969), .Q(\REGISTERS[21][6] )
         );
  DLH_X1 \REGISTERS_reg[21][5]  ( .G(n4862), .D(n4965), .Q(\REGISTERS[21][5] )
         );
  DLH_X1 \REGISTERS_reg[21][4]  ( .G(n4862), .D(n4961), .Q(\REGISTERS[21][4] )
         );
  DLH_X1 \REGISTERS_reg[21][3]  ( .G(n4862), .D(n4956), .Q(\REGISTERS[21][3] )
         );
  DLH_X1 \REGISTERS_reg[21][2]  ( .G(n4862), .D(n4952), .Q(\REGISTERS[21][2] )
         );
  DLH_X1 \REGISTERS_reg[21][1]  ( .G(n4862), .D(n4948), .Q(\REGISTERS[21][1] )
         );
  DLH_X1 \REGISTERS_reg[21][0]  ( .G(n4862), .D(n4946), .Q(\REGISTERS[21][0] )
         );
  DLH_X1 \REGISTERS_reg[22][31]  ( .G(n4859), .D(n5074), .Q(
        \REGISTERS[22][31] ) );
  DLH_X1 \REGISTERS_reg[22][30]  ( .G(n4859), .D(n5064), .Q(
        \REGISTERS[22][30] ) );
  DLH_X1 \REGISTERS_reg[22][29]  ( .G(n4857), .D(n5060), .Q(
        \REGISTERS[22][29] ) );
  DLH_X1 \REGISTERS_reg[22][28]  ( .G(n4857), .D(n5056), .Q(
        \REGISTERS[22][28] ) );
  DLH_X1 \REGISTERS_reg[22][27]  ( .G(n4857), .D(n5052), .Q(
        \REGISTERS[22][27] ) );
  DLH_X1 \REGISTERS_reg[22][26]  ( .G(n4857), .D(n5048), .Q(
        \REGISTERS[22][26] ) );
  DLH_X1 \REGISTERS_reg[22][25]  ( .G(n4857), .D(n5044), .Q(
        \REGISTERS[22][25] ) );
  DLH_X1 \REGISTERS_reg[22][24]  ( .G(n4857), .D(n5040), .Q(
        \REGISTERS[22][24] ) );
  DLH_X1 \REGISTERS_reg[22][23]  ( .G(n4857), .D(n5036), .Q(
        \REGISTERS[22][23] ) );
  DLH_X1 \REGISTERS_reg[22][22]  ( .G(n4857), .D(n5032), .Q(
        \REGISTERS[22][22] ) );
  DLH_X1 \REGISTERS_reg[22][21]  ( .G(n4857), .D(n5028), .Q(
        \REGISTERS[22][21] ) );
  DLH_X1 \REGISTERS_reg[22][20]  ( .G(n4857), .D(n5024), .Q(
        \REGISTERS[22][20] ) );
  DLH_X1 \REGISTERS_reg[22][19]  ( .G(n4856), .D(n5020), .Q(
        \REGISTERS[22][19] ) );
  DLH_X1 \REGISTERS_reg[22][18]  ( .G(n4856), .D(n5016), .Q(
        \REGISTERS[22][18] ) );
  DLH_X1 \REGISTERS_reg[22][17]  ( .G(n4856), .D(n5012), .Q(
        \REGISTERS[22][17] ) );
  DLH_X1 \REGISTERS_reg[22][16]  ( .G(n4856), .D(n5009), .Q(
        \REGISTERS[22][16] ) );
  DLH_X1 \REGISTERS_reg[22][15]  ( .G(n4856), .D(n5004), .Q(
        \REGISTERS[22][15] ) );
  DLH_X1 \REGISTERS_reg[22][14]  ( .G(n4856), .D(n5000), .Q(
        \REGISTERS[22][14] ) );
  DLH_X1 \REGISTERS_reg[22][13]  ( .G(n4856), .D(n4996), .Q(
        \REGISTERS[22][13] ) );
  DLH_X1 \REGISTERS_reg[22][12]  ( .G(n4856), .D(n4992), .Q(
        \REGISTERS[22][12] ) );
  DLH_X1 \REGISTERS_reg[22][11]  ( .G(n4856), .D(n4988), .Q(
        \REGISTERS[22][11] ) );
  DLH_X1 \REGISTERS_reg[22][10]  ( .G(n4856), .D(n4985), .Q(
        \REGISTERS[22][10] ) );
  DLH_X1 \REGISTERS_reg[22][9]  ( .G(n4858), .D(n4981), .Q(\REGISTERS[22][9] )
         );
  DLH_X1 \REGISTERS_reg[22][8]  ( .G(n4858), .D(n4976), .Q(\REGISTERS[22][8] )
         );
  DLH_X1 \REGISTERS_reg[22][7]  ( .G(n4858), .D(n4973), .Q(\REGISTERS[22][7] )
         );
  DLH_X1 \REGISTERS_reg[22][6]  ( .G(n4858), .D(n4968), .Q(\REGISTERS[22][6] )
         );
  DLH_X1 \REGISTERS_reg[22][5]  ( .G(n4858), .D(n4964), .Q(\REGISTERS[22][5] )
         );
  DLH_X1 \REGISTERS_reg[22][4]  ( .G(n4858), .D(n4960), .Q(\REGISTERS[22][4] )
         );
  DLH_X1 \REGISTERS_reg[22][3]  ( .G(n4858), .D(n4956), .Q(\REGISTERS[22][3] )
         );
  DLH_X1 \REGISTERS_reg[22][2]  ( .G(n4858), .D(n4952), .Q(\REGISTERS[22][2] )
         );
  DLH_X1 \REGISTERS_reg[22][1]  ( .G(n4858), .D(n4948), .Q(\REGISTERS[22][1] )
         );
  DLH_X1 \REGISTERS_reg[22][0]  ( .G(n4858), .D(n4944), .Q(\REGISTERS[22][0] )
         );
  DLH_X1 \REGISTERS_reg[23][31]  ( .G(n4855), .D(n5074), .Q(
        \REGISTERS[23][31] ) );
  DLH_X1 \REGISTERS_reg[23][30]  ( .G(n4855), .D(n5064), .Q(
        \REGISTERS[23][30] ) );
  DLH_X1 \REGISTERS_reg[23][29]  ( .G(n4853), .D(n5060), .Q(
        \REGISTERS[23][29] ) );
  DLH_X1 \REGISTERS_reg[23][28]  ( .G(n4853), .D(n5056), .Q(
        \REGISTERS[23][28] ) );
  DLH_X1 \REGISTERS_reg[23][27]  ( .G(n4853), .D(n5055), .Q(
        \REGISTERS[23][27] ) );
  DLH_X1 \REGISTERS_reg[23][26]  ( .G(n4853), .D(n5048), .Q(
        \REGISTERS[23][26] ) );
  DLH_X1 \REGISTERS_reg[23][25]  ( .G(n4853), .D(n5044), .Q(
        \REGISTERS[23][25] ) );
  DLH_X1 \REGISTERS_reg[23][24]  ( .G(n4853), .D(n5043), .Q(
        \REGISTERS[23][24] ) );
  DLH_X1 \REGISTERS_reg[23][23]  ( .G(n4853), .D(n5039), .Q(
        \REGISTERS[23][23] ) );
  DLH_X1 \REGISTERS_reg[23][22]  ( .G(n4853), .D(n5032), .Q(
        \REGISTERS[23][22] ) );
  DLH_X1 \REGISTERS_reg[23][21]  ( .G(n4853), .D(n5030), .Q(
        \REGISTERS[23][21] ) );
  DLH_X1 \REGISTERS_reg[23][20]  ( .G(n4853), .D(n5024), .Q(
        \REGISTERS[23][20] ) );
  DLH_X1 \REGISTERS_reg[23][19]  ( .G(n4852), .D(n5020), .Q(
        \REGISTERS[23][19] ) );
  DLH_X1 \REGISTERS_reg[23][18]  ( .G(n4852), .D(n5018), .Q(
        \REGISTERS[23][18] ) );
  DLH_X1 \REGISTERS_reg[23][17]  ( .G(n4852), .D(n5014), .Q(
        \REGISTERS[23][17] ) );
  DLH_X1 \REGISTERS_reg[23][16]  ( .G(n4852), .D(n5008), .Q(
        \REGISTERS[23][16] ) );
  DLH_X1 \REGISTERS_reg[23][15]  ( .G(n4852), .D(n5004), .Q(
        \REGISTERS[23][15] ) );
  DLH_X1 \REGISTERS_reg[23][14]  ( .G(n4852), .D(n5002), .Q(
        \REGISTERS[23][14] ) );
  DLH_X1 \REGISTERS_reg[23][13]  ( .G(n4852), .D(n4999), .Q(
        \REGISTERS[23][13] ) );
  DLH_X1 \REGISTERS_reg[23][12]  ( .G(n4852), .D(n4994), .Q(
        \REGISTERS[23][12] ) );
  DLH_X1 \REGISTERS_reg[23][11]  ( .G(n4852), .D(n4988), .Q(
        \REGISTERS[23][11] ) );
  DLH_X1 \REGISTERS_reg[23][10]  ( .G(n4852), .D(n4984), .Q(
        \REGISTERS[23][10] ) );
  DLH_X1 \REGISTERS_reg[23][9]  ( .G(n4854), .D(n4980), .Q(\REGISTERS[23][9] )
         );
  DLH_X1 \REGISTERS_reg[23][8]  ( .G(n4854), .D(n4978), .Q(\REGISTERS[23][8] )
         );
  DLH_X1 \REGISTERS_reg[23][7]  ( .G(n4854), .D(n4974), .Q(\REGISTERS[23][7] )
         );
  DLH_X1 \REGISTERS_reg[23][6]  ( .G(n4854), .D(n4970), .Q(\REGISTERS[23][6] )
         );
  DLH_X1 \REGISTERS_reg[23][5]  ( .G(n4854), .D(n4966), .Q(\REGISTERS[23][5] )
         );
  DLH_X1 \REGISTERS_reg[23][4]  ( .G(n4854), .D(n4962), .Q(\REGISTERS[23][4] )
         );
  DLH_X1 \REGISTERS_reg[23][3]  ( .G(n4854), .D(n4958), .Q(\REGISTERS[23][3] )
         );
  DLH_X1 \REGISTERS_reg[23][2]  ( .G(n4854), .D(n4954), .Q(\REGISTERS[23][2] )
         );
  DLH_X1 \REGISTERS_reg[23][1]  ( .G(n4854), .D(n4951), .Q(\REGISTERS[23][1] )
         );
  DLH_X1 \REGISTERS_reg[23][0]  ( .G(n4854), .D(n4947), .Q(\REGISTERS[23][0] )
         );
  DLH_X1 \REGISTERS_reg[24][31]  ( .G(n4851), .D(n5073), .Q(
        \REGISTERS[24][31] ) );
  DLH_X1 \REGISTERS_reg[24][30]  ( .G(n4851), .D(n5066), .Q(
        \REGISTERS[24][30] ) );
  DLH_X1 \REGISTERS_reg[24][29]  ( .G(n4849), .D(n5062), .Q(
        \REGISTERS[24][29] ) );
  DLH_X1 \REGISTERS_reg[24][28]  ( .G(n4849), .D(n5058), .Q(
        \REGISTERS[24][28] ) );
  DLH_X1 \REGISTERS_reg[24][27]  ( .G(n4849), .D(n5054), .Q(
        \REGISTERS[24][27] ) );
  DLH_X1 \REGISTERS_reg[24][26]  ( .G(n4849), .D(n5050), .Q(
        \REGISTERS[24][26] ) );
  DLH_X1 \REGISTERS_reg[24][25]  ( .G(n4849), .D(n5046), .Q(
        \REGISTERS[24][25] ) );
  DLH_X1 \REGISTERS_reg[24][24]  ( .G(n4849), .D(n5041), .Q(
        \REGISTERS[24][24] ) );
  DLH_X1 \REGISTERS_reg[24][23]  ( .G(n4849), .D(n5038), .Q(
        \REGISTERS[24][23] ) );
  DLH_X1 \REGISTERS_reg[24][22]  ( .G(n4849), .D(n5034), .Q(
        \REGISTERS[24][22] ) );
  DLH_X1 \REGISTERS_reg[24][21]  ( .G(n4849), .D(n5030), .Q(
        \REGISTERS[24][21] ) );
  DLH_X1 \REGISTERS_reg[24][20]  ( .G(n4849), .D(n5026), .Q(
        \REGISTERS[24][20] ) );
  DLH_X1 \REGISTERS_reg[24][19]  ( .G(n4848), .D(n5022), .Q(
        \REGISTERS[24][19] ) );
  DLH_X1 \REGISTERS_reg[24][18]  ( .G(n4848), .D(n5018), .Q(
        \REGISTERS[24][18] ) );
  DLH_X1 \REGISTERS_reg[24][17]  ( .G(n4848), .D(n5014), .Q(
        \REGISTERS[24][17] ) );
  DLH_X1 \REGISTERS_reg[24][16]  ( .G(n4848), .D(n5010), .Q(
        \REGISTERS[24][16] ) );
  DLH_X1 \REGISTERS_reg[24][15]  ( .G(n4848), .D(n5006), .Q(
        \REGISTERS[24][15] ) );
  DLH_X1 \REGISTERS_reg[24][14]  ( .G(n4848), .D(n5002), .Q(
        \REGISTERS[24][14] ) );
  DLH_X1 \REGISTERS_reg[24][13]  ( .G(n4848), .D(n4998), .Q(
        \REGISTERS[24][13] ) );
  DLH_X1 \REGISTERS_reg[24][12]  ( .G(n4848), .D(n4994), .Q(
        \REGISTERS[24][12] ) );
  DLH_X1 \REGISTERS_reg[24][11]  ( .G(n4848), .D(n4990), .Q(
        \REGISTERS[24][11] ) );
  DLH_X1 \REGISTERS_reg[24][10]  ( .G(n4848), .D(n4986), .Q(
        \REGISTERS[24][10] ) );
  DLH_X1 \REGISTERS_reg[24][9]  ( .G(n4850), .D(n4982), .Q(\REGISTERS[24][9] )
         );
  DLH_X1 \REGISTERS_reg[24][8]  ( .G(n4850), .D(n4978), .Q(\REGISTERS[24][8] )
         );
  DLH_X1 \REGISTERS_reg[24][7]  ( .G(n4850), .D(n4974), .Q(\REGISTERS[24][7] )
         );
  DLH_X1 \REGISTERS_reg[24][6]  ( .G(n4850), .D(n4970), .Q(\REGISTERS[24][6] )
         );
  DLH_X1 \REGISTERS_reg[24][5]  ( .G(n4850), .D(n4966), .Q(\REGISTERS[24][5] )
         );
  DLH_X1 \REGISTERS_reg[24][4]  ( .G(n4850), .D(n4960), .Q(\REGISTERS[24][4] )
         );
  DLH_X1 \REGISTERS_reg[24][3]  ( .G(n4850), .D(n4958), .Q(\REGISTERS[24][3] )
         );
  DLH_X1 \REGISTERS_reg[24][2]  ( .G(n4850), .D(n4954), .Q(\REGISTERS[24][2] )
         );
  DLH_X1 \REGISTERS_reg[24][1]  ( .G(n4850), .D(n4950), .Q(\REGISTERS[24][1] )
         );
  DLH_X1 \REGISTERS_reg[24][0]  ( .G(n4850), .D(n4946), .Q(\REGISTERS[24][0] )
         );
  DLH_X1 \REGISTERS_reg[25][31]  ( .G(n4847), .D(n5073), .Q(
        \REGISTERS[25][31] ) );
  DLH_X1 \REGISTERS_reg[25][30]  ( .G(n4847), .D(n5065), .Q(
        \REGISTERS[25][30] ) );
  DLH_X1 \REGISTERS_reg[25][29]  ( .G(n4845), .D(n5061), .Q(
        \REGISTERS[25][29] ) );
  DLH_X1 \REGISTERS_reg[25][28]  ( .G(n4845), .D(n5057), .Q(
        \REGISTERS[25][28] ) );
  DLH_X1 \REGISTERS_reg[25][27]  ( .G(n4845), .D(n5053), .Q(
        \REGISTERS[25][27] ) );
  DLH_X1 \REGISTERS_reg[25][26]  ( .G(n4845), .D(n5049), .Q(
        \REGISTERS[25][26] ) );
  DLH_X1 \REGISTERS_reg[25][25]  ( .G(n4845), .D(n5045), .Q(
        \REGISTERS[25][25] ) );
  DLH_X1 \REGISTERS_reg[25][24]  ( .G(n4845), .D(n5041), .Q(
        \REGISTERS[25][24] ) );
  DLH_X1 \REGISTERS_reg[25][23]  ( .G(n4845), .D(n5037), .Q(
        \REGISTERS[25][23] ) );
  DLH_X1 \REGISTERS_reg[25][22]  ( .G(n4845), .D(n5033), .Q(
        \REGISTERS[25][22] ) );
  DLH_X1 \REGISTERS_reg[25][21]  ( .G(n4845), .D(n5029), .Q(
        \REGISTERS[25][21] ) );
  DLH_X1 \REGISTERS_reg[25][20]  ( .G(n4845), .D(n5025), .Q(
        \REGISTERS[25][20] ) );
  DLH_X1 \REGISTERS_reg[25][19]  ( .G(n4844), .D(n5021), .Q(
        \REGISTERS[25][19] ) );
  DLH_X1 \REGISTERS_reg[25][18]  ( .G(n4844), .D(n5017), .Q(
        \REGISTERS[25][18] ) );
  DLH_X1 \REGISTERS_reg[25][17]  ( .G(n4844), .D(n5013), .Q(
        \REGISTERS[25][17] ) );
  DLH_X1 \REGISTERS_reg[25][16]  ( .G(n4844), .D(n5008), .Q(
        \REGISTERS[25][16] ) );
  DLH_X1 \REGISTERS_reg[25][15]  ( .G(n4844), .D(n5005), .Q(
        \REGISTERS[25][15] ) );
  DLH_X1 \REGISTERS_reg[25][14]  ( .G(n4844), .D(n5001), .Q(
        \REGISTERS[25][14] ) );
  DLH_X1 \REGISTERS_reg[25][13]  ( .G(n4844), .D(n4997), .Q(
        \REGISTERS[25][13] ) );
  DLH_X1 \REGISTERS_reg[25][12]  ( .G(n4844), .D(n4993), .Q(
        \REGISTERS[25][12] ) );
  DLH_X1 \REGISTERS_reg[25][11]  ( .G(n4844), .D(n4989), .Q(
        \REGISTERS[25][11] ) );
  DLH_X1 \REGISTERS_reg[25][10]  ( .G(n4844), .D(n4984), .Q(
        \REGISTERS[25][10] ) );
  DLH_X1 \REGISTERS_reg[25][9]  ( .G(n4846), .D(n4980), .Q(\REGISTERS[25][9] )
         );
  DLH_X1 \REGISTERS_reg[25][8]  ( .G(n4846), .D(n4977), .Q(\REGISTERS[25][8] )
         );
  DLH_X1 \REGISTERS_reg[25][7]  ( .G(n4846), .D(n4972), .Q(\REGISTERS[25][7] )
         );
  DLH_X1 \REGISTERS_reg[25][6]  ( .G(n4846), .D(n4969), .Q(\REGISTERS[25][6] )
         );
  DLH_X1 \REGISTERS_reg[25][5]  ( .G(n4846), .D(n4965), .Q(\REGISTERS[25][5] )
         );
  DLH_X1 \REGISTERS_reg[25][4]  ( .G(n4846), .D(n4960), .Q(\REGISTERS[25][4] )
         );
  DLH_X1 \REGISTERS_reg[25][3]  ( .G(n4846), .D(n4957), .Q(\REGISTERS[25][3] )
         );
  DLH_X1 \REGISTERS_reg[25][2]  ( .G(n4846), .D(n4953), .Q(\REGISTERS[25][2] )
         );
  DLH_X1 \REGISTERS_reg[25][1]  ( .G(n4846), .D(n4949), .Q(\REGISTERS[25][1] )
         );
  DLH_X1 \REGISTERS_reg[25][0]  ( .G(n4846), .D(n4945), .Q(\REGISTERS[25][0] )
         );
  DLH_X1 \REGISTERS_reg[26][31]  ( .G(n4843), .D(n5074), .Q(
        \REGISTERS[26][31] ) );
  DLH_X1 \REGISTERS_reg[26][30]  ( .G(n4843), .D(n5066), .Q(
        \REGISTERS[26][30] ) );
  DLH_X1 \REGISTERS_reg[26][29]  ( .G(n4841), .D(n5062), .Q(
        \REGISTERS[26][29] ) );
  DLH_X1 \REGISTERS_reg[26][28]  ( .G(n4841), .D(n5058), .Q(
        \REGISTERS[26][28] ) );
  DLH_X1 \REGISTERS_reg[26][27]  ( .G(n4841), .D(n5054), .Q(
        \REGISTERS[26][27] ) );
  DLH_X1 \REGISTERS_reg[26][26]  ( .G(n4841), .D(n5050), .Q(
        \REGISTERS[26][26] ) );
  DLH_X1 \REGISTERS_reg[26][25]  ( .G(n4841), .D(n5046), .Q(
        \REGISTERS[26][25] ) );
  DLH_X1 \REGISTERS_reg[26][24]  ( .G(n4841), .D(n5042), .Q(
        \REGISTERS[26][24] ) );
  DLH_X1 \REGISTERS_reg[26][23]  ( .G(n4841), .D(n5038), .Q(
        \REGISTERS[26][23] ) );
  DLH_X1 \REGISTERS_reg[26][22]  ( .G(n4841), .D(n5034), .Q(
        \REGISTERS[26][22] ) );
  DLH_X1 \REGISTERS_reg[26][21]  ( .G(n4841), .D(n5030), .Q(
        \REGISTERS[26][21] ) );
  DLH_X1 \REGISTERS_reg[26][20]  ( .G(n4841), .D(n5026), .Q(
        \REGISTERS[26][20] ) );
  DLH_X1 \REGISTERS_reg[26][19]  ( .G(n4840), .D(n5022), .Q(
        \REGISTERS[26][19] ) );
  DLH_X1 \REGISTERS_reg[26][18]  ( .G(n4840), .D(n5018), .Q(
        \REGISTERS[26][18] ) );
  DLH_X1 \REGISTERS_reg[26][17]  ( .G(n4840), .D(n5014), .Q(
        \REGISTERS[26][17] ) );
  DLH_X1 \REGISTERS_reg[26][16]  ( .G(n4840), .D(n5010), .Q(
        \REGISTERS[26][16] ) );
  DLH_X1 \REGISTERS_reg[26][15]  ( .G(n4840), .D(n5006), .Q(
        \REGISTERS[26][15] ) );
  DLH_X1 \REGISTERS_reg[26][14]  ( .G(n4840), .D(n5002), .Q(
        \REGISTERS[26][14] ) );
  DLH_X1 \REGISTERS_reg[26][13]  ( .G(n4840), .D(n4998), .Q(
        \REGISTERS[26][13] ) );
  DLH_X1 \REGISTERS_reg[26][12]  ( .G(n4840), .D(n4994), .Q(
        \REGISTERS[26][12] ) );
  DLH_X1 \REGISTERS_reg[26][11]  ( .G(n4840), .D(n4990), .Q(
        \REGISTERS[26][11] ) );
  DLH_X1 \REGISTERS_reg[26][10]  ( .G(n4840), .D(n4986), .Q(
        \REGISTERS[26][10] ) );
  DLH_X1 \REGISTERS_reg[26][9]  ( .G(n4842), .D(n4982), .Q(\REGISTERS[26][9] )
         );
  DLH_X1 \REGISTERS_reg[26][8]  ( .G(n4842), .D(n4978), .Q(\REGISTERS[26][8] )
         );
  DLH_X1 \REGISTERS_reg[26][7]  ( .G(n4842), .D(n4974), .Q(\REGISTERS[26][7] )
         );
  DLH_X1 \REGISTERS_reg[26][6]  ( .G(n4842), .D(n4970), .Q(\REGISTERS[26][6] )
         );
  DLH_X1 \REGISTERS_reg[26][5]  ( .G(n4842), .D(n4966), .Q(\REGISTERS[26][5] )
         );
  DLH_X1 \REGISTERS_reg[26][4]  ( .G(n4842), .D(n4962), .Q(\REGISTERS[26][4] )
         );
  DLH_X1 \REGISTERS_reg[26][3]  ( .G(n4842), .D(n4958), .Q(\REGISTERS[26][3] )
         );
  DLH_X1 \REGISTERS_reg[26][2]  ( .G(n4842), .D(n4954), .Q(\REGISTERS[26][2] )
         );
  DLH_X1 \REGISTERS_reg[26][1]  ( .G(n4842), .D(n4950), .Q(\REGISTERS[26][1] )
         );
  DLH_X1 \REGISTERS_reg[26][0]  ( .G(n4842), .D(n4946), .Q(\REGISTERS[26][0] )
         );
  DLH_X1 \REGISTERS_reg[27][31]  ( .G(n4839), .D(n5073), .Q(
        \REGISTERS[27][31] ) );
  DLH_X1 \REGISTERS_reg[27][30]  ( .G(n4839), .D(n5065), .Q(
        \REGISTERS[27][30] ) );
  DLH_X1 \REGISTERS_reg[27][29]  ( .G(n4837), .D(n5061), .Q(
        \REGISTERS[27][29] ) );
  DLH_X1 \REGISTERS_reg[27][28]  ( .G(n4837), .D(n5057), .Q(
        \REGISTERS[27][28] ) );
  DLH_X1 \REGISTERS_reg[27][27]  ( .G(n4837), .D(n5053), .Q(
        \REGISTERS[27][27] ) );
  DLH_X1 \REGISTERS_reg[27][26]  ( .G(n4837), .D(n5049), .Q(
        \REGISTERS[27][26] ) );
  DLH_X1 \REGISTERS_reg[27][25]  ( .G(n4837), .D(n5045), .Q(
        \REGISTERS[27][25] ) );
  DLH_X1 \REGISTERS_reg[27][24]  ( .G(n4837), .D(n5041), .Q(
        \REGISTERS[27][24] ) );
  DLH_X1 \REGISTERS_reg[27][23]  ( .G(n4837), .D(n5037), .Q(
        \REGISTERS[27][23] ) );
  DLH_X1 \REGISTERS_reg[27][22]  ( .G(n4837), .D(n5033), .Q(
        \REGISTERS[27][22] ) );
  DLH_X1 \REGISTERS_reg[27][21]  ( .G(n4837), .D(n5029), .Q(
        \REGISTERS[27][21] ) );
  DLH_X1 \REGISTERS_reg[27][20]  ( .G(n4837), .D(n5025), .Q(
        \REGISTERS[27][20] ) );
  DLH_X1 \REGISTERS_reg[27][19]  ( .G(n4836), .D(n5021), .Q(
        \REGISTERS[27][19] ) );
  DLH_X1 \REGISTERS_reg[27][18]  ( .G(n4836), .D(n5017), .Q(
        \REGISTERS[27][18] ) );
  DLH_X1 \REGISTERS_reg[27][17]  ( .G(n4836), .D(n5013), .Q(
        \REGISTERS[27][17] ) );
  DLH_X1 \REGISTERS_reg[27][16]  ( .G(n4836), .D(n5009), .Q(
        \REGISTERS[27][16] ) );
  DLH_X1 \REGISTERS_reg[27][15]  ( .G(n4836), .D(n5005), .Q(
        \REGISTERS[27][15] ) );
  DLH_X1 \REGISTERS_reg[27][14]  ( .G(n4836), .D(n5001), .Q(
        \REGISTERS[27][14] ) );
  DLH_X1 \REGISTERS_reg[27][13]  ( .G(n4836), .D(n4997), .Q(
        \REGISTERS[27][13] ) );
  DLH_X1 \REGISTERS_reg[27][12]  ( .G(n4836), .D(n4993), .Q(
        \REGISTERS[27][12] ) );
  DLH_X1 \REGISTERS_reg[27][11]  ( .G(n4836), .D(n4989), .Q(
        \REGISTERS[27][11] ) );
  DLH_X1 \REGISTERS_reg[27][10]  ( .G(n4836), .D(n4985), .Q(
        \REGISTERS[27][10] ) );
  DLH_X1 \REGISTERS_reg[27][9]  ( .G(n4838), .D(n4981), .Q(\REGISTERS[27][9] )
         );
  DLH_X1 \REGISTERS_reg[27][8]  ( .G(n4838), .D(n4977), .Q(\REGISTERS[27][8] )
         );
  DLH_X1 \REGISTERS_reg[27][7]  ( .G(n4838), .D(n4972), .Q(\REGISTERS[27][7] )
         );
  DLH_X1 \REGISTERS_reg[27][6]  ( .G(n4838), .D(n4969), .Q(\REGISTERS[27][6] )
         );
  DLH_X1 \REGISTERS_reg[27][5]  ( .G(n4838), .D(n4965), .Q(\REGISTERS[27][5] )
         );
  DLH_X1 \REGISTERS_reg[27][4]  ( .G(n4838), .D(n4960), .Q(\REGISTERS[27][4] )
         );
  DLH_X1 \REGISTERS_reg[27][3]  ( .G(n4838), .D(n4957), .Q(\REGISTERS[27][3] )
         );
  DLH_X1 \REGISTERS_reg[27][2]  ( .G(n4838), .D(n4953), .Q(\REGISTERS[27][2] )
         );
  DLH_X1 \REGISTERS_reg[27][1]  ( .G(n4838), .D(n4949), .Q(\REGISTERS[27][1] )
         );
  DLH_X1 \REGISTERS_reg[27][0]  ( .G(n4838), .D(n4945), .Q(\REGISTERS[27][0] )
         );
  DLH_X1 \REGISTERS_reg[28][31]  ( .G(n4835), .D(n5073), .Q(
        \REGISTERS[28][31] ) );
  DLH_X1 \REGISTERS_reg[28][30]  ( .G(n4835), .D(n5065), .Q(
        \REGISTERS[28][30] ) );
  DLH_X1 \REGISTERS_reg[28][29]  ( .G(n4833), .D(n5061), .Q(
        \REGISTERS[28][29] ) );
  DLH_X1 \REGISTERS_reg[28][28]  ( .G(n4833), .D(n5058), .Q(
        \REGISTERS[28][28] ) );
  DLH_X1 \REGISTERS_reg[28][27]  ( .G(n4833), .D(n5054), .Q(
        \REGISTERS[28][27] ) );
  DLH_X1 \REGISTERS_reg[28][26]  ( .G(n4833), .D(n5049), .Q(
        \REGISTERS[28][26] ) );
  DLH_X1 \REGISTERS_reg[28][25]  ( .G(n4833), .D(n5046), .Q(
        \REGISTERS[28][25] ) );
  DLH_X1 \REGISTERS_reg[28][24]  ( .G(n4833), .D(n5042), .Q(
        \REGISTERS[28][24] ) );
  DLH_X1 \REGISTERS_reg[28][23]  ( .G(n4833), .D(n5038), .Q(
        \REGISTERS[28][23] ) );
  DLH_X1 \REGISTERS_reg[28][22]  ( .G(n4833), .D(n5034), .Q(
        \REGISTERS[28][22] ) );
  DLH_X1 \REGISTERS_reg[28][21]  ( .G(n4833), .D(n5028), .Q(
        \REGISTERS[28][21] ) );
  DLH_X1 \REGISTERS_reg[28][20]  ( .G(n4833), .D(n5026), .Q(
        \REGISTERS[28][20] ) );
  DLH_X1 \REGISTERS_reg[28][19]  ( .G(n4832), .D(n5022), .Q(
        \REGISTERS[28][19] ) );
  DLH_X1 \REGISTERS_reg[28][18]  ( .G(n4832), .D(n5016), .Q(
        \REGISTERS[28][18] ) );
  DLH_X1 \REGISTERS_reg[28][17]  ( .G(n4832), .D(n5012), .Q(
        \REGISTERS[28][17] ) );
  DLH_X1 \REGISTERS_reg[28][16]  ( .G(n4832), .D(n5010), .Q(
        \REGISTERS[28][16] ) );
  DLH_X1 \REGISTERS_reg[28][15]  ( .G(n4832), .D(n5006), .Q(
        \REGISTERS[28][15] ) );
  DLH_X1 \REGISTERS_reg[28][14]  ( .G(n4832), .D(n5000), .Q(
        \REGISTERS[28][14] ) );
  DLH_X1 \REGISTERS_reg[28][13]  ( .G(n4832), .D(n4996), .Q(
        \REGISTERS[28][13] ) );
  DLH_X1 \REGISTERS_reg[28][12]  ( .G(n4832), .D(n4992), .Q(
        \REGISTERS[28][12] ) );
  DLH_X1 \REGISTERS_reg[28][11]  ( .G(n4832), .D(n4990), .Q(
        \REGISTERS[28][11] ) );
  DLH_X1 \REGISTERS_reg[28][10]  ( .G(n4832), .D(n4986), .Q(
        \REGISTERS[28][10] ) );
  DLH_X1 \REGISTERS_reg[28][9]  ( .G(n4834), .D(n4982), .Q(\REGISTERS[28][9] )
         );
  DLH_X1 \REGISTERS_reg[28][8]  ( .G(n4834), .D(n4976), .Q(\REGISTERS[28][8] )
         );
  DLH_X1 \REGISTERS_reg[28][7]  ( .G(n4834), .D(n4974), .Q(\REGISTERS[28][7] )
         );
  DLH_X1 \REGISTERS_reg[28][6]  ( .G(n4834), .D(n4968), .Q(\REGISTERS[28][6] )
         );
  DLH_X1 \REGISTERS_reg[28][5]  ( .G(n4834), .D(n4964), .Q(\REGISTERS[28][5] )
         );
  DLH_X1 \REGISTERS_reg[28][4]  ( .G(n4834), .D(n4961), .Q(\REGISTERS[28][4] )
         );
  DLH_X1 \REGISTERS_reg[28][3]  ( .G(n4834), .D(n4956), .Q(\REGISTERS[28][3] )
         );
  DLH_X1 \REGISTERS_reg[28][2]  ( .G(n4834), .D(n4952), .Q(\REGISTERS[28][2] )
         );
  DLH_X1 \REGISTERS_reg[28][1]  ( .G(n4834), .D(n4948), .Q(\REGISTERS[28][1] )
         );
  DLH_X1 \REGISTERS_reg[28][0]  ( .G(n4834), .D(n4944), .Q(\REGISTERS[28][0] )
         );
  DLH_X1 \REGISTERS_reg[29][31]  ( .G(n4831), .D(n5073), .Q(
        \REGISTERS[29][31] ) );
  DLH_X1 \REGISTERS_reg[29][30]  ( .G(n4831), .D(n5065), .Q(
        \REGISTERS[29][30] ) );
  DLH_X1 \REGISTERS_reg[29][29]  ( .G(n4829), .D(n5061), .Q(
        \REGISTERS[29][29] ) );
  DLH_X1 \REGISTERS_reg[29][28]  ( .G(n4829), .D(n5057), .Q(
        \REGISTERS[29][28] ) );
  DLH_X1 \REGISTERS_reg[29][27]  ( .G(n4829), .D(n5053), .Q(
        \REGISTERS[29][27] ) );
  DLH_X1 \REGISTERS_reg[29][26]  ( .G(n4829), .D(n5049), .Q(
        \REGISTERS[29][26] ) );
  DLH_X1 \REGISTERS_reg[29][25]  ( .G(n4829), .D(n5045), .Q(
        \REGISTERS[29][25] ) );
  DLH_X1 \REGISTERS_reg[29][24]  ( .G(n4829), .D(n5041), .Q(
        \REGISTERS[29][24] ) );
  DLH_X1 \REGISTERS_reg[29][23]  ( .G(n4829), .D(n5037), .Q(
        \REGISTERS[29][23] ) );
  DLH_X1 \REGISTERS_reg[29][22]  ( .G(n4829), .D(n5033), .Q(
        \REGISTERS[29][22] ) );
  DLH_X1 \REGISTERS_reg[29][21]  ( .G(n4829), .D(n5028), .Q(
        \REGISTERS[29][21] ) );
  DLH_X1 \REGISTERS_reg[29][20]  ( .G(n4829), .D(n5025), .Q(
        \REGISTERS[29][20] ) );
  DLH_X1 \REGISTERS_reg[29][19]  ( .G(n4828), .D(n5021), .Q(
        \REGISTERS[29][19] ) );
  DLH_X1 \REGISTERS_reg[29][18]  ( .G(n4828), .D(n5016), .Q(
        \REGISTERS[29][18] ) );
  DLH_X1 \REGISTERS_reg[29][17]  ( .G(n4828), .D(n5012), .Q(
        \REGISTERS[29][17] ) );
  DLH_X1 \REGISTERS_reg[29][16]  ( .G(n4828), .D(n5008), .Q(
        \REGISTERS[29][16] ) );
  DLH_X1 \REGISTERS_reg[29][15]  ( .G(n4828), .D(n5005), .Q(
        \REGISTERS[29][15] ) );
  DLH_X1 \REGISTERS_reg[29][14]  ( .G(n4828), .D(n5000), .Q(
        \REGISTERS[29][14] ) );
  DLH_X1 \REGISTERS_reg[29][13]  ( .G(n4828), .D(n4997), .Q(
        \REGISTERS[29][13] ) );
  DLH_X1 \REGISTERS_reg[29][12]  ( .G(n4828), .D(n4992), .Q(
        \REGISTERS[29][12] ) );
  DLH_X1 \REGISTERS_reg[29][11]  ( .G(n4828), .D(n4989), .Q(
        \REGISTERS[29][11] ) );
  DLH_X1 \REGISTERS_reg[29][10]  ( .G(n4828), .D(n4984), .Q(
        \REGISTERS[29][10] ) );
  DLH_X1 \REGISTERS_reg[29][9]  ( .G(n4830), .D(n4980), .Q(\REGISTERS[29][9] )
         );
  DLH_X1 \REGISTERS_reg[29][8]  ( .G(n4830), .D(n4976), .Q(\REGISTERS[29][8] )
         );
  DLH_X1 \REGISTERS_reg[29][7]  ( .G(n4830), .D(n4973), .Q(\REGISTERS[29][7] )
         );
  DLH_X1 \REGISTERS_reg[29][6]  ( .G(n4830), .D(n4968), .Q(\REGISTERS[29][6] )
         );
  DLH_X1 \REGISTERS_reg[29][5]  ( .G(n4830), .D(n4964), .Q(\REGISTERS[29][5] )
         );
  DLH_X1 \REGISTERS_reg[29][4]  ( .G(n4830), .D(n4961), .Q(\REGISTERS[29][4] )
         );
  DLH_X1 \REGISTERS_reg[29][3]  ( .G(n4830), .D(n4956), .Q(\REGISTERS[29][3] )
         );
  DLH_X1 \REGISTERS_reg[29][2]  ( .G(n4830), .D(n4952), .Q(\REGISTERS[29][2] )
         );
  DLH_X1 \REGISTERS_reg[29][1]  ( .G(n4830), .D(n4949), .Q(\REGISTERS[29][1] )
         );
  DLH_X1 \REGISTERS_reg[29][0]  ( .G(n4830), .D(n4945), .Q(\REGISTERS[29][0] )
         );
  DLH_X1 \REGISTERS_reg[30][31]  ( .G(n4827), .D(n5073), .Q(
        \REGISTERS[30][31] ) );
  DLH_X1 \REGISTERS_reg[30][30]  ( .G(n4827), .D(n5065), .Q(
        \REGISTERS[30][30] ) );
  DLH_X1 \REGISTERS_reg[30][29]  ( .G(n4825), .D(n5061), .Q(
        \REGISTERS[30][29] ) );
  DLH_X1 \REGISTERS_reg[30][28]  ( .G(n4825), .D(n5057), .Q(
        \REGISTERS[30][28] ) );
  DLH_X1 \REGISTERS_reg[30][27]  ( .G(n4825), .D(n5053), .Q(
        \REGISTERS[30][27] ) );
  DLH_X1 \REGISTERS_reg[30][26]  ( .G(n4825), .D(n5049), .Q(
        \REGISTERS[30][26] ) );
  DLH_X1 \REGISTERS_reg[30][25]  ( .G(n4825), .D(n5045), .Q(
        \REGISTERS[30][25] ) );
  DLH_X1 \REGISTERS_reg[30][24]  ( .G(n4825), .D(n5041), .Q(
        \REGISTERS[30][24] ) );
  DLH_X1 \REGISTERS_reg[30][23]  ( .G(n4825), .D(n5037), .Q(
        \REGISTERS[30][23] ) );
  DLH_X1 \REGISTERS_reg[30][22]  ( .G(n4825), .D(n5033), .Q(
        \REGISTERS[30][22] ) );
  DLH_X1 \REGISTERS_reg[30][21]  ( .G(n4825), .D(n5029), .Q(
        \REGISTERS[30][21] ) );
  DLH_X1 \REGISTERS_reg[30][20]  ( .G(n4825), .D(n5025), .Q(
        \REGISTERS[30][20] ) );
  DLH_X1 \REGISTERS_reg[30][19]  ( .G(n4824), .D(n5020), .Q(
        \REGISTERS[30][19] ) );
  DLH_X1 \REGISTERS_reg[30][18]  ( .G(n4824), .D(n5017), .Q(
        \REGISTERS[30][18] ) );
  DLH_X1 \REGISTERS_reg[30][17]  ( .G(n4824), .D(n5012), .Q(
        \REGISTERS[30][17] ) );
  DLH_X1 \REGISTERS_reg[30][16]  ( .G(n4824), .D(n5008), .Q(
        \REGISTERS[30][16] ) );
  DLH_X1 \REGISTERS_reg[30][15]  ( .G(n4824), .D(n5005), .Q(
        \REGISTERS[30][15] ) );
  DLH_X1 \REGISTERS_reg[30][14]  ( .G(n4824), .D(n5001), .Q(
        \REGISTERS[30][14] ) );
  DLH_X1 \REGISTERS_reg[30][13]  ( .G(n4824), .D(n4997), .Q(
        \REGISTERS[30][13] ) );
  DLH_X1 \REGISTERS_reg[30][12]  ( .G(n4824), .D(n4992), .Q(
        \REGISTERS[30][12] ) );
  DLH_X1 \REGISTERS_reg[30][11]  ( .G(n4824), .D(n4989), .Q(
        \REGISTERS[30][11] ) );
  DLH_X1 \REGISTERS_reg[30][10]  ( .G(n4824), .D(n4984), .Q(
        \REGISTERS[30][10] ) );
  DLH_X1 \REGISTERS_reg[30][9]  ( .G(n4826), .D(n4980), .Q(\REGISTERS[30][9] )
         );
  DLH_X1 \REGISTERS_reg[30][8]  ( .G(n4826), .D(n4976), .Q(\REGISTERS[30][8] )
         );
  DLH_X1 \REGISTERS_reg[30][7]  ( .G(n4826), .D(n4974), .Q(\REGISTERS[30][7] )
         );
  DLH_X1 \REGISTERS_reg[30][6]  ( .G(n4826), .D(n4968), .Q(\REGISTERS[30][6] )
         );
  DLH_X1 \REGISTERS_reg[30][5]  ( .G(n4826), .D(n4964), .Q(\REGISTERS[30][5] )
         );
  DLH_X1 \REGISTERS_reg[30][4]  ( .G(n4826), .D(n4961), .Q(\REGISTERS[30][4] )
         );
  DLH_X1 \REGISTERS_reg[30][3]  ( .G(n4826), .D(n4957), .Q(\REGISTERS[30][3] )
         );
  DLH_X1 \REGISTERS_reg[30][2]  ( .G(n4826), .D(n4953), .Q(\REGISTERS[30][2] )
         );
  DLH_X1 \REGISTERS_reg[30][1]  ( .G(n4826), .D(n4949), .Q(\REGISTERS[30][1] )
         );
  DLH_X1 \REGISTERS_reg[30][0]  ( .G(n4826), .D(n4944), .Q(\REGISTERS[30][0] )
         );
  DLH_X1 \REGISTERS_reg[31][31]  ( .G(n4823), .D(n5072), .Q(
        \REGISTERS[31][31] ) );
  DLH_X1 \REGISTERS_reg[31][30]  ( .G(n4823), .D(n5066), .Q(
        \REGISTERS[31][30] ) );
  DLH_X1 \REGISTERS_reg[31][29]  ( .G(n4821), .D(n5062), .Q(
        \REGISTERS[31][29] ) );
  DLH_X1 \REGISTERS_reg[31][28]  ( .G(n4821), .D(n5057), .Q(
        \REGISTERS[31][28] ) );
  DLH_X1 \REGISTERS_reg[31][27]  ( .G(n4821), .D(n5053), .Q(
        \REGISTERS[31][27] ) );
  DLH_X1 \REGISTERS_reg[31][26]  ( .G(n4821), .D(n5050), .Q(
        \REGISTERS[31][26] ) );
  DLH_X1 \REGISTERS_reg[31][25]  ( .G(n4821), .D(n5045), .Q(
        \REGISTERS[31][25] ) );
  DLH_X1 \REGISTERS_reg[31][24]  ( .G(n4821), .D(n5040), .Q(
        \REGISTERS[31][24] ) );
  DLH_X1 \REGISTERS_reg[31][23]  ( .G(n4821), .D(n5037), .Q(
        \REGISTERS[31][23] ) );
  DLH_X1 \REGISTERS_reg[31][22]  ( .G(n4821), .D(n5033), .Q(
        \REGISTERS[31][22] ) );
  DLH_X1 \REGISTERS_reg[31][21]  ( .G(n4821), .D(n5030), .Q(
        \REGISTERS[31][21] ) );
  DLH_X1 \REGISTERS_reg[31][20]  ( .G(n4821), .D(n5025), .Q(
        \REGISTERS[31][20] ) );
  DLH_X1 \REGISTERS_reg[31][19]  ( .G(n4820), .D(n5020), .Q(
        \REGISTERS[31][19] ) );
  DLH_X1 \REGISTERS_reg[31][18]  ( .G(n4820), .D(n5018), .Q(
        \REGISTERS[31][18] ) );
  DLH_X1 \REGISTERS_reg[31][17]  ( .G(n4820), .D(n5014), .Q(
        \REGISTERS[31][17] ) );
  DLH_X1 \REGISTERS_reg[31][16]  ( .G(n4820), .D(n5010), .Q(
        \REGISTERS[31][16] ) );
  DLH_X1 \REGISTERS_reg[31][15]  ( .G(n4820), .D(n5005), .Q(
        \REGISTERS[31][15] ) );
  DLH_X1 \REGISTERS_reg[31][14]  ( .G(n4820), .D(n5002), .Q(
        \REGISTERS[31][14] ) );
  DLH_X1 \REGISTERS_reg[31][13]  ( .G(n4820), .D(n4997), .Q(
        \REGISTERS[31][13] ) );
  DLH_X1 \REGISTERS_reg[31][12]  ( .G(n4820), .D(n4994), .Q(
        \REGISTERS[31][12] ) );
  DLH_X1 \REGISTERS_reg[31][11]  ( .G(n4820), .D(n4989), .Q(
        \REGISTERS[31][11] ) );
  DLH_X1 \REGISTERS_reg[31][10]  ( .G(n4820), .D(n4986), .Q(
        \REGISTERS[31][10] ) );
  DLH_X1 \REGISTERS_reg[31][9]  ( .G(n4822), .D(n4982), .Q(\REGISTERS[31][9] )
         );
  DLH_X1 \REGISTERS_reg[31][8]  ( .G(n4822), .D(n4978), .Q(\REGISTERS[31][8] )
         );
  DLH_X1 \REGISTERS_reg[31][7]  ( .G(n4822), .D(n4974), .Q(\REGISTERS[31][7] )
         );
  DLH_X1 \REGISTERS_reg[31][6]  ( .G(n4822), .D(n4970), .Q(\REGISTERS[31][6] )
         );
  DLH_X1 \REGISTERS_reg[31][5]  ( .G(n4822), .D(n4966), .Q(\REGISTERS[31][5] )
         );
  DLH_X1 \REGISTERS_reg[31][4]  ( .G(n4822), .D(n4961), .Q(\REGISTERS[31][4] )
         );
  DLH_X1 \REGISTERS_reg[31][3]  ( .G(n4822), .D(n4958), .Q(\REGISTERS[31][3] )
         );
  DLH_X1 \REGISTERS_reg[31][2]  ( .G(n4822), .D(n4954), .Q(\REGISTERS[31][2] )
         );
  DLH_X1 \REGISTERS_reg[31][1]  ( .G(n4822), .D(n4949), .Q(\REGISTERS[31][1] )
         );
  DLH_X1 \REGISTERS_reg[31][0]  ( .G(n4822), .D(n4945), .Q(\REGISTERS[31][0] )
         );
  DLH_X1 \OUT1_reg[31]  ( .G(n4815), .D(N2481), .Q(OUT1[31]) );
  DLH_X1 \OUT1_reg[30]  ( .G(n4814), .D(N2479), .Q(OUT1[30]) );
  DLH_X1 \OUT1_reg[29]  ( .G(n4812), .D(N2477), .Q(OUT1[29]) );
  DLH_X1 \OUT1_reg[28]  ( .G(n4815), .D(N2475), .Q(OUT1[28]) );
  DLH_X1 \OUT1_reg[27]  ( .G(n4814), .D(N2473), .Q(OUT1[27]) );
  DLH_X1 \OUT1_reg[26]  ( .G(n4812), .D(N2471), .Q(OUT1[26]) );
  DLH_X1 \OUT1_reg[25]  ( .G(n4812), .D(N2469), .Q(OUT1[25]) );
  DLH_X1 \OUT1_reg[24]  ( .G(n4814), .D(N2467), .Q(OUT1[24]) );
  DLH_X1 \OUT1_reg[23]  ( .G(n4813), .D(N2465), .Q(OUT1[23]) );
  DLH_X1 \OUT1_reg[22]  ( .G(n4812), .D(N2463), .Q(OUT1[22]) );
  DLH_X1 \OUT1_reg[21]  ( .G(n4812), .D(N2461), .Q(OUT1[21]) );
  DLH_X1 \OUT1_reg[20]  ( .G(n4812), .D(N2459), .Q(OUT1[20]) );
  DLH_X1 \OUT1_reg[19]  ( .G(n4812), .D(N2457), .Q(OUT1[19]) );
  DLH_X1 \OUT1_reg[18]  ( .G(n4814), .D(N2455), .Q(OUT1[18]) );
  DLH_X1 \OUT1_reg[17]  ( .G(n4814), .D(N2453), .Q(OUT1[17]) );
  DLH_X1 \OUT1_reg[16]  ( .G(n4814), .D(N2451), .Q(OUT1[16]) );
  DLH_X1 \OUT1_reg[15]  ( .G(n4814), .D(N2449), .Q(OUT1[15]) );
  DLH_X1 \OUT1_reg[14]  ( .G(n4813), .D(N2447), .Q(OUT1[14]) );
  DLH_X1 \OUT1_reg[13]  ( .G(n4813), .D(N2445), .Q(OUT1[13]) );
  DLH_X1 \OUT1_reg[12]  ( .G(n4813), .D(N2443), .Q(OUT1[12]) );
  DLH_X1 \OUT1_reg[11]  ( .G(n4812), .D(N2441), .Q(OUT1[11]) );
  DLH_X1 \OUT1_reg[10]  ( .G(n4814), .D(N2439), .Q(OUT1[10]) );
  DLH_X1 \OUT1_reg[9]  ( .G(n4813), .D(N2437), .Q(OUT1[9]) );
  DLH_X1 \OUT1_reg[8]  ( .G(n4813), .D(N2435), .Q(OUT1[8]) );
  DLH_X1 \OUT1_reg[7]  ( .G(n4813), .D(N2433), .Q(OUT1[7]) );
  DLH_X1 \OUT1_reg[6]  ( .G(n4813), .D(N2431), .Q(OUT1[6]) );
  DLH_X1 \OUT1_reg[5]  ( .G(n4812), .D(N2429), .Q(OUT1[5]) );
  DLH_X1 \OUT1_reg[4]  ( .G(n4813), .D(N2427), .Q(OUT1[4]) );
  DLH_X1 \OUT1_reg[3]  ( .G(n4814), .D(N2425), .Q(OUT1[3]) );
  DLH_X1 \OUT1_reg[2]  ( .G(n4814), .D(N2423), .Q(OUT1[2]) );
  DLH_X1 \OUT1_reg[1]  ( .G(n4813), .D(N2421), .Q(OUT1[1]) );
  DLH_X1 \OUT1_reg[0]  ( .G(n4812), .D(N2419), .Q(OUT1[0]) );
  DLH_X1 \OUT2_reg[31]  ( .G(n4817), .D(N2545), .Q(OUT2[31]) );
  DLH_X1 \OUT2_reg[30]  ( .G(n4819), .D(N2543), .Q(OUT2[30]) );
  DLH_X1 \OUT2_reg[29]  ( .G(n4818), .D(N2541), .Q(OUT2[29]) );
  DLH_X1 \OUT2_reg[28]  ( .G(n4817), .D(N2539), .Q(OUT2[28]) );
  DLH_X1 \OUT2_reg[27]  ( .G(n4817), .D(N2537), .Q(OUT2[27]) );
  DLH_X1 \OUT2_reg[26]  ( .G(n4817), .D(N2535), .Q(OUT2[26]) );
  DLH_X1 \OUT2_reg[25]  ( .G(n4817), .D(N2533), .Q(OUT2[25]) );
  DLH_X1 \OUT2_reg[24]  ( .G(n4817), .D(N2531), .Q(OUT2[24]) );
  DLH_X1 \OUT2_reg[23]  ( .G(n4818), .D(N2529), .Q(OUT2[23]) );
  DLH_X1 \OUT2_reg[22]  ( .G(n4817), .D(N2527), .Q(OUT2[22]) );
  DLH_X1 \OUT2_reg[21]  ( .G(n4816), .D(N2525), .Q(OUT2[21]) );
  DLH_X1 \OUT2_reg[20]  ( .G(n4819), .D(N2523), .Q(OUT2[20]) );
  DLH_X1 \OUT2_reg[19]  ( .G(n4816), .D(N2521), .Q(OUT2[19]) );
  DLH_X1 \OUT2_reg[18]  ( .G(n4816), .D(N2519), .Q(OUT2[18]) );
  DLH_X1 \OUT2_reg[17]  ( .G(n4816), .D(N2517), .Q(OUT2[17]) );
  DLH_X1 \OUT2_reg[16]  ( .G(n4817), .D(N2515), .Q(OUT2[16]) );
  DLH_X1 \OUT2_reg[15]  ( .G(n4816), .D(N2513), .Q(OUT2[15]) );
  DLH_X1 \OUT2_reg[14]  ( .G(n4818), .D(N2511), .Q(OUT2[14]) );
  DLH_X1 \OUT2_reg[13]  ( .G(n4816), .D(N2509), .Q(OUT2[13]) );
  DLH_X1 \OUT2_reg[12]  ( .G(n4818), .D(N2507), .Q(OUT2[12]) );
  DLH_X1 \OUT2_reg[11]  ( .G(n4816), .D(N2505), .Q(OUT2[11]) );
  DLH_X1 \OUT2_reg[10]  ( .G(n4816), .D(N2503), .Q(OUT2[10]) );
  DLH_X1 \OUT2_reg[9]  ( .G(n4818), .D(N2501), .Q(OUT2[9]) );
  DLH_X1 \OUT2_reg[8]  ( .G(n4818), .D(N2499), .Q(OUT2[8]) );
  DLH_X1 \OUT2_reg[7]  ( .G(n4818), .D(N2497), .Q(OUT2[7]) );
  DLH_X1 \OUT2_reg[6]  ( .G(n4818), .D(N2495), .Q(OUT2[6]) );
  DLH_X1 \OUT2_reg[5]  ( .G(n4818), .D(N2493), .Q(OUT2[5]) );
  DLH_X1 \OUT2_reg[4]  ( .G(n4816), .D(N2491), .Q(OUT2[4]) );
  DLH_X1 \OUT2_reg[3]  ( .G(n4817), .D(N2489), .Q(OUT2[3]) );
  DLH_X1 \OUT2_reg[2]  ( .G(n4817), .D(N2487), .Q(OUT2[2]) );
  DLH_X1 \OUT2_reg[1]  ( .G(n4818), .D(N2485), .Q(OUT2[1]) );
  DLH_X1 \OUT2_reg[0]  ( .G(n4816), .D(N2483), .Q(OUT2[0]) );
  NOR3_X2 U727 ( .A1(n525), .A2(ADD_RD2[2]), .A3(n1676), .ZN(n1647) );
  NOR3_X2 U1894 ( .A1(n525), .A2(ADD_RD1[2]), .A3(n2301), .ZN(n2283) );
  NAND3_X1 U1899 ( .A1(ADD_WR[3]), .A2(n535), .A3(ADD_WR[4]), .ZN(n526) );
  NAND3_X1 U1900 ( .A1(n535), .A2(n537), .A3(ADD_WR[4]), .ZN(n536) );
  NAND3_X1 U1901 ( .A1(n535), .A2(n539), .A3(ADD_WR[3]), .ZN(n538) );
  NAND3_X1 U1902 ( .A1(ADD_WR[1]), .A2(ADD_WR[0]), .A3(ADD_WR[2]), .ZN(n527)
         );
  NAND3_X1 U1903 ( .A1(ADD_WR[1]), .A2(n541), .A3(ADD_WR[2]), .ZN(n528) );
  NAND3_X1 U1904 ( .A1(ADD_WR[0]), .A2(n542), .A3(ADD_WR[2]), .ZN(n529) );
  NAND3_X1 U1905 ( .A1(n541), .A2(n542), .A3(ADD_WR[2]), .ZN(n530) );
  NAND3_X1 U1906 ( .A1(ADD_WR[0]), .A2(n543), .A3(ADD_WR[1]), .ZN(n531) );
  NAND3_X1 U1907 ( .A1(n541), .A2(n543), .A3(ADD_WR[1]), .ZN(n532) );
  NAND3_X1 U1908 ( .A1(n542), .A2(n543), .A3(ADD_WR[0]), .ZN(n533) );
  NAND3_X1 U1909 ( .A1(n537), .A2(n539), .A3(n535), .ZN(n540) );
  NAND3_X1 U1910 ( .A1(n542), .A2(n543), .A3(n541), .ZN(n534) );
  NOR3_X1 U3 ( .A1(ADD_RD2[1]), .A2(ADD_RD2[2]), .A3(n525), .ZN(n1646) );
  NOR3_X1 U4 ( .A1(ADD_RD1[1]), .A2(ADD_RD1[2]), .A3(n525), .ZN(n2282) );
  BUF_X1 U5 ( .A(n5076), .Z(n5080) );
  BUF_X1 U6 ( .A(n5077), .Z(n5081) );
  BUF_X1 U7 ( .A(n5076), .Z(n5079) );
  BUF_X1 U8 ( .A(n5076), .Z(n5078) );
  BUF_X1 U9 ( .A(n5077), .Z(n5082) );
  BUF_X1 U10 ( .A(RESET), .Z(n5076) );
  BUF_X1 U11 ( .A(RESET), .Z(n5077) );
  BUF_X1 U12 ( .A(n1689), .Z(n4707) );
  BUF_X1 U13 ( .A(n1694), .Z(n4695) );
  BUF_X1 U14 ( .A(n1699), .Z(n4683) );
  BUF_X1 U15 ( .A(n1704), .Z(n4671) );
  BUF_X1 U16 ( .A(n1713), .Z(n4659) );
  BUF_X1 U17 ( .A(n1718), .Z(n4647) );
  BUF_X1 U18 ( .A(n1723), .Z(n4635) );
  BUF_X1 U19 ( .A(n1728), .Z(n4623) );
  BUF_X1 U20 ( .A(n1689), .Z(n4708) );
  BUF_X1 U21 ( .A(n1694), .Z(n4696) );
  BUF_X1 U22 ( .A(n1699), .Z(n4684) );
  BUF_X1 U23 ( .A(n1704), .Z(n4672) );
  BUF_X1 U24 ( .A(n1713), .Z(n4660) );
  BUF_X1 U25 ( .A(n1718), .Z(n4648) );
  BUF_X1 U26 ( .A(n1723), .Z(n4636) );
  BUF_X1 U27 ( .A(n1728), .Z(n4624) );
  BUF_X1 U28 ( .A(n1686), .Z(n4713) );
  BUF_X1 U29 ( .A(n1691), .Z(n4701) );
  BUF_X1 U30 ( .A(n1696), .Z(n4689) );
  BUF_X1 U31 ( .A(n1701), .Z(n4677) );
  BUF_X1 U32 ( .A(n1710), .Z(n4665) );
  BUF_X1 U33 ( .A(n1715), .Z(n4653) );
  BUF_X1 U34 ( .A(n1720), .Z(n4641) );
  BUF_X1 U35 ( .A(n1725), .Z(n4629) );
  BUF_X1 U36 ( .A(n552), .Z(n4806) );
  BUF_X1 U37 ( .A(n559), .Z(n4794) );
  BUF_X1 U38 ( .A(n605), .Z(n4722) );
  BUF_X1 U39 ( .A(n566), .Z(n4782) );
  BUF_X1 U40 ( .A(n573), .Z(n4770) );
  BUF_X1 U41 ( .A(n584), .Z(n4758) );
  BUF_X1 U42 ( .A(n591), .Z(n4746) );
  BUF_X1 U43 ( .A(n598), .Z(n4734) );
  BUF_X1 U44 ( .A(n552), .Z(n4807) );
  BUF_X1 U45 ( .A(n559), .Z(n4795) );
  BUF_X1 U46 ( .A(n566), .Z(n4783) );
  BUF_X1 U47 ( .A(n573), .Z(n4771) );
  BUF_X1 U48 ( .A(n584), .Z(n4759) );
  BUF_X1 U49 ( .A(n591), .Z(n4747) );
  BUF_X1 U50 ( .A(n598), .Z(n4735) );
  BUF_X1 U51 ( .A(n605), .Z(n4723) );
  BUF_X1 U52 ( .A(n1690), .Z(n4704) );
  BUF_X1 U53 ( .A(n1695), .Z(n4692) );
  BUF_X1 U54 ( .A(n1700), .Z(n4680) );
  BUF_X1 U55 ( .A(n1705), .Z(n4668) );
  BUF_X1 U56 ( .A(n1714), .Z(n4656) );
  BUF_X1 U57 ( .A(n1719), .Z(n4644) );
  BUF_X1 U58 ( .A(n1724), .Z(n4632) );
  BUF_X1 U59 ( .A(n1729), .Z(n4620) );
  BUF_X1 U60 ( .A(n1690), .Z(n4705) );
  BUF_X1 U61 ( .A(n1695), .Z(n4693) );
  BUF_X1 U62 ( .A(n1700), .Z(n4681) );
  BUF_X1 U63 ( .A(n1705), .Z(n4669) );
  BUF_X1 U64 ( .A(n1714), .Z(n4657) );
  BUF_X1 U65 ( .A(n1719), .Z(n4645) );
  BUF_X1 U66 ( .A(n1724), .Z(n4633) );
  BUF_X1 U67 ( .A(n1729), .Z(n4621) );
  OAI21_X1 U68 ( .B1(n526), .B2(n527), .A(n5079), .ZN(n4604) );
  OAI21_X1 U69 ( .B1(n526), .B2(n528), .A(n5078), .ZN(n4600) );
  OAI21_X1 U70 ( .B1(n526), .B2(n529), .A(n5078), .ZN(n4596) );
  OAI21_X1 U71 ( .B1(n526), .B2(n530), .A(n5078), .ZN(n4592) );
  OAI21_X1 U72 ( .B1(n526), .B2(n531), .A(n5078), .ZN(n4588) );
  OAI21_X1 U73 ( .B1(n526), .B2(n532), .A(n5078), .ZN(n4584) );
  OAI21_X1 U74 ( .B1(n526), .B2(n533), .A(n5078), .ZN(n4580) );
  OAI21_X1 U75 ( .B1(n526), .B2(n534), .A(n5078), .ZN(n4576) );
  BUF_X1 U76 ( .A(n1692), .Z(n4700) );
  BUF_X1 U77 ( .A(n1716), .Z(n4652) );
  BUF_X1 U78 ( .A(n1726), .Z(n4628) );
  BUF_X1 U79 ( .A(n1687), .Z(n4712) );
  BUF_X1 U80 ( .A(n1697), .Z(n4688) );
  BUF_X1 U81 ( .A(n1702), .Z(n4676) );
  BUF_X1 U82 ( .A(n1711), .Z(n4664) );
  BUF_X1 U83 ( .A(n1721), .Z(n4640) );
  BUF_X1 U84 ( .A(n1689), .Z(n4709) );
  BUF_X1 U85 ( .A(n1694), .Z(n4697) );
  BUF_X1 U86 ( .A(n1704), .Z(n4673) );
  BUF_X1 U87 ( .A(n1699), .Z(n4685) );
  BUF_X1 U88 ( .A(n1713), .Z(n4661) );
  BUF_X1 U89 ( .A(n1718), .Z(n4649) );
  BUF_X1 U90 ( .A(n1723), .Z(n4637) );
  BUF_X1 U91 ( .A(n1728), .Z(n4625) );
  BUF_X1 U92 ( .A(n1686), .Z(n4715) );
  BUF_X1 U93 ( .A(n1691), .Z(n4703) );
  BUF_X1 U94 ( .A(n1696), .Z(n4691) );
  BUF_X1 U95 ( .A(n1701), .Z(n4679) );
  BUF_X1 U96 ( .A(n1710), .Z(n4667) );
  BUF_X1 U97 ( .A(n1715), .Z(n4655) );
  BUF_X1 U98 ( .A(n1720), .Z(n4643) );
  BUF_X1 U99 ( .A(n1725), .Z(n4631) );
  BUF_X1 U100 ( .A(n557), .Z(n4797) );
  BUF_X1 U101 ( .A(n589), .Z(n4749) );
  BUF_X1 U102 ( .A(n603), .Z(n4725) );
  BUF_X1 U103 ( .A(n557), .Z(n4798) );
  BUF_X1 U104 ( .A(n589), .Z(n4750) );
  BUF_X1 U105 ( .A(n603), .Z(n4726) );
  BUF_X1 U106 ( .A(n555), .Z(n4803) );
  BUF_X1 U107 ( .A(n562), .Z(n4791) );
  BUF_X1 U108 ( .A(n569), .Z(n4779) );
  BUF_X1 U109 ( .A(n576), .Z(n4767) );
  BUF_X1 U110 ( .A(n587), .Z(n4755) );
  BUF_X1 U111 ( .A(n594), .Z(n4743) );
  BUF_X1 U112 ( .A(n601), .Z(n4731) );
  BUF_X1 U113 ( .A(n608), .Z(n4719) );
  BUF_X1 U114 ( .A(n555), .Z(n4804) );
  BUF_X1 U115 ( .A(n562), .Z(n4792) );
  BUF_X1 U116 ( .A(n569), .Z(n4780) );
  BUF_X1 U117 ( .A(n576), .Z(n4768) );
  BUF_X1 U118 ( .A(n587), .Z(n4756) );
  BUF_X1 U119 ( .A(n594), .Z(n4744) );
  BUF_X1 U120 ( .A(n601), .Z(n4732) );
  BUF_X1 U121 ( .A(n608), .Z(n4720) );
  BUF_X1 U122 ( .A(n550), .Z(n4809) );
  BUF_X1 U123 ( .A(n564), .Z(n4785) );
  BUF_X1 U124 ( .A(n571), .Z(n4773) );
  BUF_X1 U125 ( .A(n582), .Z(n4761) );
  BUF_X1 U126 ( .A(n596), .Z(n4737) );
  BUF_X1 U127 ( .A(n550), .Z(n4810) );
  BUF_X1 U128 ( .A(n564), .Z(n4786) );
  BUF_X1 U129 ( .A(n571), .Z(n4774) );
  BUF_X1 U130 ( .A(n582), .Z(n4762) );
  BUF_X1 U131 ( .A(n596), .Z(n4738) );
  BUF_X1 U132 ( .A(n556), .Z(n4800) );
  BUF_X1 U133 ( .A(n563), .Z(n4788) );
  BUF_X1 U134 ( .A(n570), .Z(n4776) );
  BUF_X1 U135 ( .A(n577), .Z(n4764) );
  BUF_X1 U136 ( .A(n588), .Z(n4752) );
  BUF_X1 U137 ( .A(n595), .Z(n4740) );
  BUF_X1 U138 ( .A(n602), .Z(n4728) );
  BUF_X1 U139 ( .A(n609), .Z(n4716) );
  BUF_X1 U140 ( .A(n556), .Z(n4801) );
  BUF_X1 U141 ( .A(n563), .Z(n4789) );
  BUF_X1 U142 ( .A(n570), .Z(n4777) );
  BUF_X1 U143 ( .A(n577), .Z(n4765) );
  BUF_X1 U144 ( .A(n588), .Z(n4753) );
  BUF_X1 U145 ( .A(n595), .Z(n4741) );
  BUF_X1 U146 ( .A(n602), .Z(n4729) );
  BUF_X1 U147 ( .A(n609), .Z(n4717) );
  BUF_X1 U148 ( .A(n559), .Z(n4796) );
  BUF_X1 U149 ( .A(n591), .Z(n4748) );
  BUF_X1 U150 ( .A(n552), .Z(n4808) );
  BUF_X1 U151 ( .A(n573), .Z(n4772) );
  BUF_X1 U152 ( .A(n566), .Z(n4784) );
  BUF_X1 U153 ( .A(n584), .Z(n4760) );
  BUF_X1 U154 ( .A(n598), .Z(n4736) );
  BUF_X1 U155 ( .A(n605), .Z(n4724) );
  BUF_X1 U156 ( .A(n1690), .Z(n4706) );
  BUF_X1 U157 ( .A(n1695), .Z(n4694) );
  BUF_X1 U158 ( .A(n1700), .Z(n4682) );
  BUF_X1 U159 ( .A(n1705), .Z(n4670) );
  BUF_X1 U160 ( .A(n1714), .Z(n4658) );
  BUF_X1 U161 ( .A(n1719), .Z(n4646) );
  BUF_X1 U162 ( .A(n1724), .Z(n4634) );
  BUF_X1 U163 ( .A(n1729), .Z(n4622) );
  OAI21_X1 U164 ( .B1(n527), .B2(n536), .A(n5078), .ZN(n4572) );
  OAI21_X1 U165 ( .B1(n528), .B2(n536), .A(n5078), .ZN(n4568) );
  OAI21_X1 U166 ( .B1(n529), .B2(n536), .A(n5079), .ZN(n4564) );
  OAI21_X1 U167 ( .B1(n530), .B2(n536), .A(n5078), .ZN(n4560) );
  OAI21_X1 U168 ( .B1(n531), .B2(n536), .A(n5079), .ZN(n4556) );
  OAI21_X1 U169 ( .B1(n532), .B2(n536), .A(n5079), .ZN(n4552) );
  OAI21_X1 U170 ( .B1(n533), .B2(n536), .A(n5079), .ZN(n4548) );
  OAI21_X1 U171 ( .B1(n534), .B2(n536), .A(n5079), .ZN(n4544) );
  OAI21_X1 U172 ( .B1(n527), .B2(n538), .A(n5079), .ZN(n4540) );
  OAI21_X1 U173 ( .B1(n528), .B2(n538), .A(n5079), .ZN(n4536) );
  OAI21_X1 U174 ( .B1(n529), .B2(n538), .A(n5079), .ZN(n4532) );
  OAI21_X1 U175 ( .B1(n530), .B2(n538), .A(n5079), .ZN(n4528) );
  OAI21_X1 U176 ( .B1(n531), .B2(n538), .A(n5079), .ZN(n4524) );
  OAI21_X1 U177 ( .B1(n532), .B2(n538), .A(n5080), .ZN(n4520) );
  OAI21_X1 U178 ( .B1(n533), .B2(n538), .A(n5080), .ZN(n4516) );
  OAI21_X1 U179 ( .B1(n534), .B2(n538), .A(n5080), .ZN(n4512) );
  OAI21_X1 U180 ( .B1(n527), .B2(n540), .A(n5080), .ZN(n4508) );
  OAI21_X1 U181 ( .B1(n528), .B2(n540), .A(n5080), .ZN(n4504) );
  OAI21_X1 U182 ( .B1(n529), .B2(n540), .A(n5080), .ZN(n4500) );
  OAI21_X1 U183 ( .B1(n530), .B2(n540), .A(n5080), .ZN(n4496) );
  OAI21_X1 U184 ( .B1(n531), .B2(n540), .A(n5080), .ZN(n4492) );
  OAI21_X1 U185 ( .B1(n532), .B2(n540), .A(n5080), .ZN(n4488) );
  OAI21_X1 U186 ( .B1(n533), .B2(n540), .A(n5080), .ZN(n4484) );
  OAI21_X1 U187 ( .B1(n534), .B2(n540), .A(n5078), .ZN(n4356) );
  BUF_X1 U188 ( .A(n557), .Z(n4799) );
  BUF_X1 U189 ( .A(n589), .Z(n4751) );
  BUF_X1 U190 ( .A(n603), .Z(n4727) );
  BUF_X1 U191 ( .A(n571), .Z(n4775) );
  BUF_X1 U192 ( .A(n550), .Z(n4811) );
  BUF_X1 U193 ( .A(n555), .Z(n4805) );
  BUF_X1 U194 ( .A(n562), .Z(n4793) );
  BUF_X1 U195 ( .A(n576), .Z(n4769) );
  BUF_X1 U196 ( .A(n569), .Z(n4781) );
  BUF_X1 U197 ( .A(n587), .Z(n4757) );
  BUF_X1 U198 ( .A(n594), .Z(n4745) );
  BUF_X1 U199 ( .A(n601), .Z(n4733) );
  BUF_X1 U200 ( .A(n608), .Z(n4721) );
  BUF_X1 U201 ( .A(n564), .Z(n4787) );
  BUF_X1 U202 ( .A(n582), .Z(n4763) );
  BUF_X1 U203 ( .A(n596), .Z(n4739) );
  BUF_X1 U204 ( .A(n556), .Z(n4802) );
  BUF_X1 U205 ( .A(n563), .Z(n4790) );
  BUF_X1 U206 ( .A(n570), .Z(n4778) );
  BUF_X1 U207 ( .A(n577), .Z(n4766) );
  BUF_X1 U208 ( .A(n588), .Z(n4754) );
  BUF_X1 U209 ( .A(n595), .Z(n4742) );
  BUF_X1 U210 ( .A(n602), .Z(n4730) );
  BUF_X1 U211 ( .A(n609), .Z(n4718) );
  BUF_X1 U212 ( .A(n1692), .Z(n4698) );
  BUF_X1 U213 ( .A(n1716), .Z(n4650) );
  BUF_X1 U214 ( .A(n1726), .Z(n4626) );
  BUF_X1 U215 ( .A(n1692), .Z(n4699) );
  BUF_X1 U216 ( .A(n1716), .Z(n4651) );
  BUF_X1 U217 ( .A(n1726), .Z(n4627) );
  BUF_X1 U218 ( .A(n1687), .Z(n4710) );
  BUF_X1 U219 ( .A(n1697), .Z(n4686) );
  BUF_X1 U220 ( .A(n1702), .Z(n4674) );
  BUF_X1 U221 ( .A(n1711), .Z(n4662) );
  BUF_X1 U222 ( .A(n1721), .Z(n4638) );
  BUF_X1 U223 ( .A(n1687), .Z(n4711) );
  BUF_X1 U224 ( .A(n1697), .Z(n4687) );
  BUF_X1 U225 ( .A(n1702), .Z(n4675) );
  BUF_X1 U226 ( .A(n1711), .Z(n4663) );
  BUF_X1 U227 ( .A(n1721), .Z(n4639) );
  BUF_X1 U228 ( .A(n1686), .Z(n4714) );
  BUF_X1 U229 ( .A(n1691), .Z(n4702) );
  BUF_X1 U230 ( .A(n1696), .Z(n4690) );
  BUF_X1 U231 ( .A(n1701), .Z(n4678) );
  BUF_X1 U232 ( .A(n1710), .Z(n4666) );
  BUF_X1 U233 ( .A(n1715), .Z(n4654) );
  BUF_X1 U234 ( .A(n1720), .Z(n4642) );
  BUF_X1 U235 ( .A(n1725), .Z(n4630) );
  NAND2_X1 U236 ( .A1(n1647), .A2(n1653), .ZN(n571) );
  NAND2_X1 U237 ( .A1(n2283), .A2(n2286), .ZN(n1702) );
  NAND2_X1 U238 ( .A1(n2283), .A2(n2287), .ZN(n1701) );
  NAND2_X1 U239 ( .A1(n1647), .A2(n1652), .ZN(n573) );
  NAND2_X1 U240 ( .A1(n1641), .A2(n1647), .ZN(n557) );
  NAND2_X1 U241 ( .A1(n1666), .A2(n1647), .ZN(n589) );
  NAND2_X1 U242 ( .A1(n1674), .A2(n1647), .ZN(n603) );
  NAND2_X1 U243 ( .A1(n2277), .A2(n2283), .ZN(n1692) );
  NAND2_X1 U244 ( .A1(n2295), .A2(n2283), .ZN(n1716) );
  NAND2_X1 U245 ( .A1(n2299), .A2(n2283), .ZN(n1726) );
  NAND2_X1 U246 ( .A1(n2279), .A2(n2283), .ZN(n1691) );
  NAND2_X1 U247 ( .A1(n2296), .A2(n2283), .ZN(n1715) );
  NAND2_X1 U248 ( .A1(n2300), .A2(n2283), .ZN(n1725) );
  NAND2_X1 U249 ( .A1(n1639), .A2(n1647), .ZN(n559) );
  NAND2_X1 U250 ( .A1(n1665), .A2(n1647), .ZN(n591) );
  NAND2_X1 U251 ( .A1(n1673), .A2(n1647), .ZN(n605) );
  NAND2_X1 U252 ( .A1(n1666), .A2(n1642), .ZN(n582) );
  NAND2_X1 U253 ( .A1(n1674), .A2(n1642), .ZN(n596) );
  NAND2_X1 U254 ( .A1(n2295), .A2(n2280), .ZN(n1711) );
  NAND2_X1 U255 ( .A1(n2299), .A2(n2280), .ZN(n1721) );
  NAND2_X1 U256 ( .A1(n2296), .A2(n2280), .ZN(n1710) );
  NAND2_X1 U257 ( .A1(n2300), .A2(n2280), .ZN(n1720) );
  NAND2_X1 U258 ( .A1(n1642), .A2(n1653), .ZN(n564) );
  NAND2_X1 U259 ( .A1(n2280), .A2(n2286), .ZN(n1697) );
  NAND2_X1 U260 ( .A1(n1665), .A2(n1642), .ZN(n584) );
  NAND2_X1 U261 ( .A1(n1673), .A2(n1642), .ZN(n598) );
  NAND2_X1 U262 ( .A1(n1641), .A2(n1642), .ZN(n550) );
  NAND2_X1 U263 ( .A1(n2277), .A2(n2280), .ZN(n1687) );
  NAND2_X1 U264 ( .A1(n2280), .A2(n2287), .ZN(n1696) );
  AND2_X1 U265 ( .A1(n1646), .A2(n1653), .ZN(n576) );
  BUF_X1 U266 ( .A(n4436), .Z(n4989) );
  BUF_X1 U267 ( .A(n4388), .Z(n5037) );
  BUF_X1 U268 ( .A(n4372), .Z(n5053) );
  BUF_X1 U269 ( .A(n4464), .Z(n4962) );
  BUF_X1 U270 ( .A(n4472), .Z(n4954) );
  BUF_X1 U271 ( .A(n4468), .Z(n4958) );
  BUF_X1 U272 ( .A(n4444), .Z(n4982) );
  BUF_X1 U273 ( .A(n4440), .Z(n4986) );
  BUF_X1 U274 ( .A(n4424), .Z(n5002) );
  BUF_X1 U275 ( .A(n4416), .Z(n5010) );
  BUF_X1 U276 ( .A(n4408), .Z(n5018) );
  BUF_X1 U277 ( .A(n4396), .Z(n5030) );
  BUF_X1 U278 ( .A(n4352), .Z(n5074) );
  BUF_X1 U279 ( .A(n4404), .Z(n5021) );
  BUF_X1 U280 ( .A(n4376), .Z(n5050) );
  BUF_X1 U281 ( .A(n4364), .Z(n5062) );
  BUF_X1 U282 ( .A(n4360), .Z(n5066) );
  BUF_X1 U283 ( .A(n4480), .Z(n4944) );
  BUF_X1 U284 ( .A(n4460), .Z(n4964) );
  BUF_X1 U285 ( .A(n4456), .Z(n4968) );
  BUF_X1 U286 ( .A(n4448), .Z(n4976) );
  BUF_X1 U287 ( .A(n4432), .Z(n4992) );
  BUF_X1 U288 ( .A(n4412), .Z(n5012) );
  BUF_X1 U289 ( .A(n4400), .Z(n5026) );
  BUF_X1 U290 ( .A(n4392), .Z(n5034) );
  BUF_X1 U291 ( .A(n4384), .Z(n5041) );
  BUF_X1 U292 ( .A(n4380), .Z(n5046) );
  BUF_X1 U293 ( .A(n4368), .Z(n5058) );
  BUF_X1 U294 ( .A(n4476), .Z(n4949) );
  BUF_X1 U295 ( .A(n4472), .Z(n4953) );
  BUF_X1 U296 ( .A(n4468), .Z(n4957) );
  BUF_X1 U297 ( .A(n4452), .Z(n4973) );
  BUF_X1 U298 ( .A(n4428), .Z(n4997) );
  BUF_X1 U299 ( .A(n4424), .Z(n5001) );
  BUF_X1 U300 ( .A(n4420), .Z(n5006) );
  BUF_X1 U301 ( .A(n4408), .Z(n5017) );
  BUF_X1 U302 ( .A(n4400), .Z(n5025) );
  BUF_X1 U303 ( .A(n4396), .Z(n5029) );
  BUF_X1 U304 ( .A(n4392), .Z(n5033) );
  BUF_X1 U305 ( .A(n4380), .Z(n5045) );
  BUF_X1 U306 ( .A(n4368), .Z(n5057) );
  BUF_X1 U307 ( .A(n4476), .Z(n4948) );
  BUF_X1 U308 ( .A(n4472), .Z(n4952) );
  BUF_X1 U309 ( .A(n4468), .Z(n4956) );
  BUF_X1 U310 ( .A(n4464), .Z(n4961) );
  BUF_X1 U311 ( .A(n4460), .Z(n4966) );
  BUF_X1 U312 ( .A(n4456), .Z(n4970) );
  BUF_X1 U313 ( .A(n4452), .Z(n4974) );
  BUF_X1 U314 ( .A(n4448), .Z(n4978) );
  BUF_X1 U315 ( .A(n4444), .Z(n4980) );
  BUF_X1 U316 ( .A(n4440), .Z(n4984) );
  BUF_X1 U317 ( .A(n4432), .Z(n4994) );
  BUF_X1 U318 ( .A(n4428), .Z(n4996) );
  BUF_X1 U319 ( .A(n4424), .Z(n5000) );
  BUF_X1 U320 ( .A(n4420), .Z(n5004) );
  BUF_X1 U321 ( .A(n4416), .Z(n5008) );
  BUF_X1 U322 ( .A(n4412), .Z(n5014) );
  BUF_X1 U323 ( .A(n4408), .Z(n5016) );
  BUF_X1 U324 ( .A(n4396), .Z(n5028) );
  BUF_X1 U325 ( .A(n4376), .Z(n5049) );
  BUF_X1 U326 ( .A(n4364), .Z(n5061) );
  BUF_X1 U327 ( .A(n4360), .Z(n5065) );
  BUF_X1 U328 ( .A(n4352), .Z(n5073) );
  BUF_X1 U329 ( .A(n4480), .Z(n4945) );
  BUF_X1 U330 ( .A(n4460), .Z(n4965) );
  BUF_X1 U331 ( .A(n4456), .Z(n4969) );
  BUF_X1 U332 ( .A(n4448), .Z(n4977) );
  BUF_X1 U333 ( .A(n4444), .Z(n4981) );
  BUF_X1 U334 ( .A(n4440), .Z(n4985) );
  BUF_X1 U335 ( .A(n4436), .Z(n4988) );
  BUF_X1 U336 ( .A(n4432), .Z(n4993) );
  BUF_X1 U337 ( .A(n4416), .Z(n5009) );
  BUF_X1 U338 ( .A(n4412), .Z(n5013) );
  BUF_X1 U339 ( .A(n4404), .Z(n5020) );
  BUF_X1 U340 ( .A(n4388), .Z(n5036) );
  BUF_X1 U341 ( .A(n4384), .Z(n5040) );
  BUF_X1 U342 ( .A(n4372), .Z(n5052) );
  BUF_X1 U343 ( .A(n4480), .Z(n4946) );
  BUF_X1 U344 ( .A(n4476), .Z(n4950) );
  BUF_X1 U345 ( .A(n4464), .Z(n4960) );
  BUF_X1 U346 ( .A(n4452), .Z(n4972) );
  BUF_X1 U347 ( .A(n4436), .Z(n4990) );
  BUF_X1 U348 ( .A(n4428), .Z(n4998) );
  BUF_X1 U349 ( .A(n4420), .Z(n5005) );
  BUF_X1 U350 ( .A(n4404), .Z(n5022) );
  BUF_X1 U351 ( .A(n4400), .Z(n5024) );
  BUF_X1 U352 ( .A(n4392), .Z(n5032) );
  BUF_X1 U353 ( .A(n4388), .Z(n5038) );
  BUF_X1 U354 ( .A(n4384), .Z(n5042) );
  BUF_X1 U355 ( .A(n4380), .Z(n5044) );
  BUF_X1 U356 ( .A(n4376), .Z(n5048) );
  BUF_X1 U357 ( .A(n4372), .Z(n5054) );
  BUF_X1 U358 ( .A(n4368), .Z(n5056) );
  BUF_X1 U359 ( .A(n4364), .Z(n5060) );
  BUF_X1 U360 ( .A(n4360), .Z(n5064) );
  BUF_X1 U361 ( .A(n4352), .Z(n5072) );
  AND2_X1 U362 ( .A1(n1641), .A2(n1646), .ZN(n562) );
  AND2_X1 U363 ( .A1(n1639), .A2(n1646), .ZN(n563) );
  AND2_X1 U364 ( .A1(n1652), .A2(n1646), .ZN(n577) );
  AND2_X1 U365 ( .A1(n1666), .A2(n1646), .ZN(n594) );
  AND2_X1 U366 ( .A1(n1665), .A2(n1646), .ZN(n595) );
  AND2_X1 U367 ( .A1(n1674), .A2(n1646), .ZN(n608) );
  AND2_X1 U368 ( .A1(n1673), .A2(n1646), .ZN(n609) );
  AND2_X1 U369 ( .A1(n1666), .A2(n1640), .ZN(n587) );
  AND2_X1 U370 ( .A1(n1665), .A2(n1640), .ZN(n588) );
  AND2_X1 U371 ( .A1(n1674), .A2(n1640), .ZN(n601) );
  AND2_X1 U372 ( .A1(n1673), .A2(n1640), .ZN(n602) );
  NAND2_X1 U373 ( .A1(n1642), .A2(n1652), .ZN(n566) );
  INV_X1 U374 ( .A(n525), .ZN(n1675) );
  AND2_X1 U375 ( .A1(n1640), .A2(n1653), .ZN(n569) );
  AND2_X1 U376 ( .A1(n1640), .A2(n1652), .ZN(n570) );
  AND2_X1 U377 ( .A1(n1641), .A2(n1640), .ZN(n555) );
  AND2_X1 U378 ( .A1(n1639), .A2(n1640), .ZN(n556) );
  NAND2_X1 U379 ( .A1(n2279), .A2(n2280), .ZN(n1686) );
  NAND2_X1 U380 ( .A1(n1639), .A2(n1642), .ZN(n552) );
  AND2_X1 U381 ( .A1(n2282), .A2(n2287), .ZN(n1704) );
  INV_X1 U382 ( .A(ADD_WR[2]), .ZN(n543) );
  INV_X1 U383 ( .A(ADD_WR[0]), .ZN(n541) );
  INV_X1 U384 ( .A(ADD_WR[1]), .ZN(n542) );
  AND2_X1 U385 ( .A1(n2279), .A2(n2282), .ZN(n1694) );
  AND2_X1 U386 ( .A1(n2277), .A2(n2282), .ZN(n1695) );
  AND2_X1 U387 ( .A1(n2286), .A2(n2282), .ZN(n1705) );
  AND2_X1 U388 ( .A1(n2296), .A2(n2282), .ZN(n1718) );
  AND2_X1 U389 ( .A1(n2295), .A2(n2282), .ZN(n1719) );
  AND2_X1 U390 ( .A1(n2300), .A2(n2282), .ZN(n1728) );
  AND2_X1 U391 ( .A1(n2299), .A2(n2282), .ZN(n1729) );
  AND2_X1 U392 ( .A1(n2296), .A2(n2278), .ZN(n1713) );
  AND2_X1 U393 ( .A1(n2295), .A2(n2278), .ZN(n1714) );
  AND2_X1 U394 ( .A1(n2300), .A2(n2278), .ZN(n1723) );
  AND2_X1 U395 ( .A1(n2299), .A2(n2278), .ZN(n1724) );
  NAND2_X1 U396 ( .A1(n1874), .A2(n1875), .ZN(N2463) );
  NOR4_X1 U397 ( .A1(n1884), .A2(n1885), .A3(n1886), .A4(n1887), .ZN(n1874) );
  NOR4_X1 U398 ( .A1(n1876), .A2(n1877), .A3(n1878), .A4(n1879), .ZN(n1875) );
  OAI221_X1 U399 ( .B1(n913), .B2(n4631), .C1(n914), .C2(n4628), .A(n1891), 
        .ZN(n1884) );
  NAND2_X1 U400 ( .A1(n1856), .A2(n1857), .ZN(N2465) );
  NOR4_X1 U401 ( .A1(n1866), .A2(n1867), .A3(n1868), .A4(n1869), .ZN(n1856) );
  NOR4_X1 U402 ( .A1(n1858), .A2(n1859), .A3(n1860), .A4(n1861), .ZN(n1857) );
  OAI221_X1 U403 ( .B1(n879), .B2(n4631), .C1(n880), .C2(n4628), .A(n1873), 
        .ZN(n1866) );
  NAND2_X1 U404 ( .A1(n1838), .A2(n1839), .ZN(N2467) );
  NOR4_X1 U405 ( .A1(n1848), .A2(n1849), .A3(n1850), .A4(n1851), .ZN(n1838) );
  NOR4_X1 U406 ( .A1(n1840), .A2(n1841), .A3(n1842), .A4(n1843), .ZN(n1839) );
  OAI221_X1 U407 ( .B1(n845), .B2(n4631), .C1(n846), .C2(n4628), .A(n1855), 
        .ZN(n1848) );
  NAND2_X1 U408 ( .A1(n1820), .A2(n1821), .ZN(N2469) );
  NOR4_X1 U409 ( .A1(n1830), .A2(n1831), .A3(n1832), .A4(n1833), .ZN(n1820) );
  NOR4_X1 U410 ( .A1(n1822), .A2(n1823), .A3(n1824), .A4(n1825), .ZN(n1821) );
  OAI221_X1 U411 ( .B1(n811), .B2(n4631), .C1(n812), .C2(n4628), .A(n1837), 
        .ZN(n1830) );
  NAND2_X1 U412 ( .A1(n1802), .A2(n1803), .ZN(N2471) );
  NOR4_X1 U413 ( .A1(n1812), .A2(n1813), .A3(n1814), .A4(n1815), .ZN(n1802) );
  NOR4_X1 U414 ( .A1(n1804), .A2(n1805), .A3(n1806), .A4(n1807), .ZN(n1803) );
  OAI221_X1 U415 ( .B1(n777), .B2(n4631), .C1(n778), .C2(n4628), .A(n1819), 
        .ZN(n1812) );
  NAND2_X1 U416 ( .A1(n1784), .A2(n1785), .ZN(N2473) );
  NOR4_X1 U417 ( .A1(n1794), .A2(n1795), .A3(n1796), .A4(n1797), .ZN(n1784) );
  NOR4_X1 U418 ( .A1(n1786), .A2(n1787), .A3(n1788), .A4(n1789), .ZN(n1785) );
  OAI221_X1 U419 ( .B1(n743), .B2(n4631), .C1(n744), .C2(n4628), .A(n1801), 
        .ZN(n1794) );
  NAND2_X1 U420 ( .A1(n1766), .A2(n1767), .ZN(N2475) );
  NOR4_X1 U421 ( .A1(n1776), .A2(n1777), .A3(n1778), .A4(n1779), .ZN(n1766) );
  NOR4_X1 U422 ( .A1(n1768), .A2(n1769), .A3(n1770), .A4(n1771), .ZN(n1767) );
  OAI221_X1 U423 ( .B1(n709), .B2(n4631), .C1(n710), .C2(n4628), .A(n1783), 
        .ZN(n1776) );
  NAND2_X1 U424 ( .A1(n1748), .A2(n1749), .ZN(N2477) );
  NOR4_X1 U425 ( .A1(n1758), .A2(n1759), .A3(n1760), .A4(n1761), .ZN(n1748) );
  NOR4_X1 U426 ( .A1(n1750), .A2(n1751), .A3(n1752), .A4(n1753), .ZN(n1749) );
  OAI221_X1 U427 ( .B1(n675), .B2(n4631), .C1(n676), .C2(n4628), .A(n1765), 
        .ZN(n1758) );
  NAND2_X1 U428 ( .A1(n1730), .A2(n1731), .ZN(N2479) );
  NOR4_X1 U429 ( .A1(n1740), .A2(n1741), .A3(n1742), .A4(n1743), .ZN(n1730) );
  NOR4_X1 U430 ( .A1(n1732), .A2(n1733), .A3(n1734), .A4(n1735), .ZN(n1731) );
  OAI221_X1 U431 ( .B1(n641), .B2(n4631), .C1(n642), .C2(n4628), .A(n1747), 
        .ZN(n1740) );
  NAND2_X1 U432 ( .A1(n1680), .A2(n1681), .ZN(N2481) );
  NOR4_X1 U433 ( .A1(n1706), .A2(n1707), .A3(n1708), .A4(n1709), .ZN(n1680) );
  NOR4_X1 U434 ( .A1(n1682), .A2(n1683), .A3(n1684), .A4(n1685), .ZN(n1681) );
  OAI221_X1 U435 ( .B1(n604), .B2(n4631), .C1(n606), .C2(n4628), .A(n1727), 
        .ZN(n1706) );
  NAND2_X1 U436 ( .A1(n2270), .A2(n2271), .ZN(N2419) );
  NOR4_X1 U437 ( .A1(n2290), .A2(n2291), .A3(n2292), .A4(n2293), .ZN(n2270) );
  NOR4_X1 U438 ( .A1(n2272), .A2(n2273), .A3(n2274), .A4(n2275), .ZN(n2271) );
  OAI221_X1 U439 ( .B1(n1677), .B2(n4629), .C1(n1678), .C2(n4626), .A(n2302), 
        .ZN(n2290) );
  NAND2_X1 U440 ( .A1(n2252), .A2(n2253), .ZN(N2421) );
  NOR4_X1 U441 ( .A1(n2262), .A2(n2263), .A3(n2264), .A4(n2265), .ZN(n2252) );
  NOR4_X1 U442 ( .A1(n2254), .A2(n2255), .A3(n2256), .A4(n2257), .ZN(n2253) );
  OAI221_X1 U443 ( .B1(n1627), .B2(n4629), .C1(n1628), .C2(n4626), .A(n2269), 
        .ZN(n2262) );
  NAND2_X1 U444 ( .A1(n2234), .A2(n2235), .ZN(N2423) );
  NOR4_X1 U445 ( .A1(n2244), .A2(n2245), .A3(n2246), .A4(n2247), .ZN(n2234) );
  NOR4_X1 U446 ( .A1(n2236), .A2(n2237), .A3(n2238), .A4(n2239), .ZN(n2235) );
  OAI221_X1 U447 ( .B1(n1593), .B2(n4629), .C1(n1594), .C2(n4626), .A(n2251), 
        .ZN(n2244) );
  NAND2_X1 U448 ( .A1(n2216), .A2(n2217), .ZN(N2425) );
  NOR4_X1 U449 ( .A1(n2226), .A2(n2227), .A3(n2228), .A4(n2229), .ZN(n2216) );
  NOR4_X1 U450 ( .A1(n2218), .A2(n2219), .A3(n2220), .A4(n2221), .ZN(n2217) );
  OAI221_X1 U451 ( .B1(n1559), .B2(n4629), .C1(n1560), .C2(n4626), .A(n2233), 
        .ZN(n2226) );
  NAND2_X1 U452 ( .A1(n2198), .A2(n2199), .ZN(N2427) );
  NOR4_X1 U453 ( .A1(n2208), .A2(n2209), .A3(n2210), .A4(n2211), .ZN(n2198) );
  NOR4_X1 U454 ( .A1(n2200), .A2(n2201), .A3(n2202), .A4(n2203), .ZN(n2199) );
  OAI221_X1 U455 ( .B1(n1525), .B2(n4629), .C1(n1526), .C2(n4626), .A(n2215), 
        .ZN(n2208) );
  NAND2_X1 U456 ( .A1(n2180), .A2(n2181), .ZN(N2429) );
  NOR4_X1 U457 ( .A1(n2190), .A2(n2191), .A3(n2192), .A4(n2193), .ZN(n2180) );
  NOR4_X1 U458 ( .A1(n2182), .A2(n2183), .A3(n2184), .A4(n2185), .ZN(n2181) );
  OAI221_X1 U459 ( .B1(n1491), .B2(n4629), .C1(n1492), .C2(n4626), .A(n2197), 
        .ZN(n2190) );
  NAND2_X1 U460 ( .A1(n2162), .A2(n2163), .ZN(N2431) );
  NOR4_X1 U461 ( .A1(n2172), .A2(n2173), .A3(n2174), .A4(n2175), .ZN(n2162) );
  NOR4_X1 U462 ( .A1(n2164), .A2(n2165), .A3(n2166), .A4(n2167), .ZN(n2163) );
  OAI221_X1 U463 ( .B1(n1457), .B2(n4629), .C1(n1458), .C2(n4626), .A(n2179), 
        .ZN(n2172) );
  NAND2_X1 U464 ( .A1(n2144), .A2(n2145), .ZN(N2433) );
  NOR4_X1 U465 ( .A1(n2154), .A2(n2155), .A3(n2156), .A4(n2157), .ZN(n2144) );
  NOR4_X1 U466 ( .A1(n2146), .A2(n2147), .A3(n2148), .A4(n2149), .ZN(n2145) );
  OAI221_X1 U467 ( .B1(n1423), .B2(n4629), .C1(n1424), .C2(n4626), .A(n2161), 
        .ZN(n2154) );
  NAND2_X1 U468 ( .A1(n2126), .A2(n2127), .ZN(N2435) );
  NOR4_X1 U469 ( .A1(n2136), .A2(n2137), .A3(n2138), .A4(n2139), .ZN(n2126) );
  NOR4_X1 U470 ( .A1(n2128), .A2(n2129), .A3(n2130), .A4(n2131), .ZN(n2127) );
  OAI221_X1 U471 ( .B1(n1389), .B2(n4629), .C1(n1390), .C2(n4626), .A(n2143), 
        .ZN(n2136) );
  NAND2_X1 U472 ( .A1(n2108), .A2(n2109), .ZN(N2437) );
  NOR4_X1 U473 ( .A1(n2118), .A2(n2119), .A3(n2120), .A4(n2121), .ZN(n2108) );
  NOR4_X1 U474 ( .A1(n2110), .A2(n2111), .A3(n2112), .A4(n2113), .ZN(n2109) );
  OAI221_X1 U475 ( .B1(n1355), .B2(n4629), .C1(n1356), .C2(n4626), .A(n2125), 
        .ZN(n2118) );
  NAND2_X1 U476 ( .A1(n2090), .A2(n2091), .ZN(N2439) );
  NOR4_X1 U477 ( .A1(n2100), .A2(n2101), .A3(n2102), .A4(n2103), .ZN(n2090) );
  NOR4_X1 U478 ( .A1(n2092), .A2(n2093), .A3(n2094), .A4(n2095), .ZN(n2091) );
  OAI221_X1 U479 ( .B1(n1321), .B2(n4629), .C1(n1322), .C2(n4626), .A(n2107), 
        .ZN(n2100) );
  NAND2_X1 U480 ( .A1(n2072), .A2(n2073), .ZN(N2441) );
  NOR4_X1 U481 ( .A1(n2082), .A2(n2083), .A3(n2084), .A4(n2085), .ZN(n2072) );
  NOR4_X1 U482 ( .A1(n2074), .A2(n2075), .A3(n2076), .A4(n2077), .ZN(n2073) );
  OAI221_X1 U483 ( .B1(n1287), .B2(n4630), .C1(n1288), .C2(n4627), .A(n2089), 
        .ZN(n2082) );
  NAND2_X1 U484 ( .A1(n2054), .A2(n2055), .ZN(N2443) );
  NOR4_X1 U485 ( .A1(n2064), .A2(n2065), .A3(n2066), .A4(n2067), .ZN(n2054) );
  NOR4_X1 U486 ( .A1(n2056), .A2(n2057), .A3(n2058), .A4(n2059), .ZN(n2055) );
  OAI221_X1 U487 ( .B1(n1253), .B2(n4630), .C1(n1254), .C2(n4627), .A(n2071), 
        .ZN(n2064) );
  NAND2_X1 U488 ( .A1(n2036), .A2(n2037), .ZN(N2445) );
  NOR4_X1 U489 ( .A1(n2046), .A2(n2047), .A3(n2048), .A4(n2049), .ZN(n2036) );
  NOR4_X1 U490 ( .A1(n2038), .A2(n2039), .A3(n2040), .A4(n2041), .ZN(n2037) );
  OAI221_X1 U491 ( .B1(n1219), .B2(n4630), .C1(n1220), .C2(n4627), .A(n2053), 
        .ZN(n2046) );
  NAND2_X1 U492 ( .A1(n2018), .A2(n2019), .ZN(N2447) );
  NOR4_X1 U493 ( .A1(n2028), .A2(n2029), .A3(n2030), .A4(n2031), .ZN(n2018) );
  NOR4_X1 U494 ( .A1(n2020), .A2(n2021), .A3(n2022), .A4(n2023), .ZN(n2019) );
  OAI221_X1 U495 ( .B1(n1185), .B2(n4630), .C1(n1186), .C2(n4627), .A(n2035), 
        .ZN(n2028) );
  NAND2_X1 U496 ( .A1(n2000), .A2(n2001), .ZN(N2449) );
  NOR4_X1 U497 ( .A1(n2010), .A2(n2011), .A3(n2012), .A4(n2013), .ZN(n2000) );
  NOR4_X1 U498 ( .A1(n2002), .A2(n2003), .A3(n2004), .A4(n2005), .ZN(n2001) );
  OAI221_X1 U499 ( .B1(n1151), .B2(n4630), .C1(n1152), .C2(n4627), .A(n2017), 
        .ZN(n2010) );
  NAND2_X1 U500 ( .A1(n1982), .A2(n1983), .ZN(N2451) );
  NOR4_X1 U501 ( .A1(n1992), .A2(n1993), .A3(n1994), .A4(n1995), .ZN(n1982) );
  NOR4_X1 U502 ( .A1(n1984), .A2(n1985), .A3(n1986), .A4(n1987), .ZN(n1983) );
  OAI221_X1 U503 ( .B1(n1117), .B2(n4630), .C1(n1118), .C2(n4627), .A(n1999), 
        .ZN(n1992) );
  NAND2_X1 U504 ( .A1(n1964), .A2(n1965), .ZN(N2453) );
  NOR4_X1 U505 ( .A1(n1974), .A2(n1975), .A3(n1976), .A4(n1977), .ZN(n1964) );
  NOR4_X1 U506 ( .A1(n1966), .A2(n1967), .A3(n1968), .A4(n1969), .ZN(n1965) );
  OAI221_X1 U507 ( .B1(n1083), .B2(n4630), .C1(n1084), .C2(n4627), .A(n1981), 
        .ZN(n1974) );
  NAND2_X1 U508 ( .A1(n1946), .A2(n1947), .ZN(N2455) );
  NOR4_X1 U509 ( .A1(n1956), .A2(n1957), .A3(n1958), .A4(n1959), .ZN(n1946) );
  NOR4_X1 U510 ( .A1(n1948), .A2(n1949), .A3(n1950), .A4(n1951), .ZN(n1947) );
  OAI221_X1 U511 ( .B1(n1049), .B2(n4630), .C1(n1050), .C2(n4627), .A(n1963), 
        .ZN(n1956) );
  NAND2_X1 U512 ( .A1(n1928), .A2(n1929), .ZN(N2457) );
  NOR4_X1 U513 ( .A1(n1938), .A2(n1939), .A3(n1940), .A4(n1941), .ZN(n1928) );
  NOR4_X1 U514 ( .A1(n1930), .A2(n1931), .A3(n1932), .A4(n1933), .ZN(n1929) );
  OAI221_X1 U515 ( .B1(n1015), .B2(n4630), .C1(n1016), .C2(n4627), .A(n1945), 
        .ZN(n1938) );
  NAND2_X1 U516 ( .A1(n1910), .A2(n1911), .ZN(N2459) );
  NOR4_X1 U517 ( .A1(n1920), .A2(n1921), .A3(n1922), .A4(n1923), .ZN(n1910) );
  NOR4_X1 U518 ( .A1(n1912), .A2(n1913), .A3(n1914), .A4(n1915), .ZN(n1911) );
  OAI221_X1 U519 ( .B1(n981), .B2(n4630), .C1(n982), .C2(n4627), .A(n1927), 
        .ZN(n1920) );
  NAND2_X1 U520 ( .A1(n1892), .A2(n1893), .ZN(N2461) );
  NOR4_X1 U521 ( .A1(n1902), .A2(n1903), .A3(n1904), .A4(n1905), .ZN(n1892) );
  NOR4_X1 U522 ( .A1(n1894), .A2(n1895), .A3(n1896), .A4(n1897), .ZN(n1893) );
  OAI221_X1 U523 ( .B1(n947), .B2(n4630), .C1(n948), .C2(n4627), .A(n1909), 
        .ZN(n1902) );
  NAND2_X1 U524 ( .A1(n1630), .A2(n1631), .ZN(N2483) );
  NOR4_X1 U525 ( .A1(n1658), .A2(n1659), .A3(n1660), .A4(n1661), .ZN(n1630) );
  NOR4_X1 U526 ( .A1(n1632), .A2(n1633), .A3(n1634), .A4(n1635), .ZN(n1631) );
  OAI221_X1 U527 ( .B1(n4725), .B2(n1677), .C1(n4722), .C2(n1678), .A(n1679), 
        .ZN(n1658) );
  NAND2_X1 U528 ( .A1(n1596), .A2(n1597), .ZN(N2485) );
  NOR4_X1 U529 ( .A1(n1614), .A2(n1615), .A3(n1616), .A4(n1617), .ZN(n1596) );
  NOR4_X1 U530 ( .A1(n1598), .A2(n1599), .A3(n1600), .A4(n1601), .ZN(n1597) );
  OAI221_X1 U531 ( .B1(n4725), .B2(n1627), .C1(n4722), .C2(n1628), .A(n1629), 
        .ZN(n1614) );
  NAND2_X1 U532 ( .A1(n1562), .A2(n1563), .ZN(N2487) );
  NOR4_X1 U533 ( .A1(n1580), .A2(n1581), .A3(n1582), .A4(n1583), .ZN(n1562) );
  NOR4_X1 U534 ( .A1(n1564), .A2(n1565), .A3(n1566), .A4(n1567), .ZN(n1563) );
  OAI221_X1 U535 ( .B1(n4725), .B2(n1593), .C1(n4722), .C2(n1594), .A(n1595), 
        .ZN(n1580) );
  NAND2_X1 U536 ( .A1(n1528), .A2(n1529), .ZN(N2489) );
  NOR4_X1 U537 ( .A1(n1546), .A2(n1547), .A3(n1548), .A4(n1549), .ZN(n1528) );
  NOR4_X1 U538 ( .A1(n1530), .A2(n1531), .A3(n1532), .A4(n1533), .ZN(n1529) );
  OAI221_X1 U539 ( .B1(n4725), .B2(n1559), .C1(n4722), .C2(n1560), .A(n1561), 
        .ZN(n1546) );
  NAND2_X1 U540 ( .A1(n1494), .A2(n1495), .ZN(N2491) );
  NOR4_X1 U541 ( .A1(n1512), .A2(n1513), .A3(n1514), .A4(n1515), .ZN(n1494) );
  NOR4_X1 U542 ( .A1(n1496), .A2(n1497), .A3(n1498), .A4(n1499), .ZN(n1495) );
  OAI221_X1 U543 ( .B1(n4725), .B2(n1525), .C1(n4722), .C2(n1526), .A(n1527), 
        .ZN(n1512) );
  NAND2_X1 U544 ( .A1(n1460), .A2(n1461), .ZN(N2493) );
  NOR4_X1 U545 ( .A1(n1478), .A2(n1479), .A3(n1480), .A4(n1481), .ZN(n1460) );
  NOR4_X1 U546 ( .A1(n1462), .A2(n1463), .A3(n1464), .A4(n1465), .ZN(n1461) );
  OAI221_X1 U547 ( .B1(n4725), .B2(n1491), .C1(n4722), .C2(n1492), .A(n1493), 
        .ZN(n1478) );
  NAND2_X1 U548 ( .A1(n1426), .A2(n1427), .ZN(N2495) );
  NOR4_X1 U549 ( .A1(n1444), .A2(n1445), .A3(n1446), .A4(n1447), .ZN(n1426) );
  NOR4_X1 U550 ( .A1(n1428), .A2(n1429), .A3(n1430), .A4(n1431), .ZN(n1427) );
  OAI221_X1 U551 ( .B1(n4725), .B2(n1457), .C1(n4722), .C2(n1458), .A(n1459), 
        .ZN(n1444) );
  NAND2_X1 U552 ( .A1(n1392), .A2(n1393), .ZN(N2497) );
  NOR4_X1 U553 ( .A1(n1410), .A2(n1411), .A3(n1412), .A4(n1413), .ZN(n1392) );
  NOR4_X1 U554 ( .A1(n1394), .A2(n1395), .A3(n1396), .A4(n1397), .ZN(n1393) );
  OAI221_X1 U555 ( .B1(n4725), .B2(n1423), .C1(n4722), .C2(n1424), .A(n1425), 
        .ZN(n1410) );
  NAND2_X1 U556 ( .A1(n1358), .A2(n1359), .ZN(N2499) );
  NOR4_X1 U557 ( .A1(n1376), .A2(n1377), .A3(n1378), .A4(n1379), .ZN(n1358) );
  NOR4_X1 U558 ( .A1(n1360), .A2(n1361), .A3(n1362), .A4(n1363), .ZN(n1359) );
  OAI221_X1 U559 ( .B1(n4725), .B2(n1389), .C1(n4722), .C2(n1390), .A(n1391), 
        .ZN(n1376) );
  NAND2_X1 U560 ( .A1(n1324), .A2(n1325), .ZN(N2501) );
  NOR4_X1 U561 ( .A1(n1342), .A2(n1343), .A3(n1344), .A4(n1345), .ZN(n1324) );
  NOR4_X1 U562 ( .A1(n1326), .A2(n1327), .A3(n1328), .A4(n1329), .ZN(n1325) );
  OAI221_X1 U563 ( .B1(n4725), .B2(n1355), .C1(n4722), .C2(n1356), .A(n1357), 
        .ZN(n1342) );
  NAND2_X1 U564 ( .A1(n1290), .A2(n1291), .ZN(N2503) );
  NOR4_X1 U565 ( .A1(n1308), .A2(n1309), .A3(n1310), .A4(n1311), .ZN(n1290) );
  NOR4_X1 U566 ( .A1(n1292), .A2(n1293), .A3(n1294), .A4(n1295), .ZN(n1291) );
  OAI221_X1 U567 ( .B1(n4725), .B2(n1321), .C1(n4722), .C2(n1322), .A(n1323), 
        .ZN(n1308) );
  NAND2_X1 U568 ( .A1(n1256), .A2(n1257), .ZN(N2505) );
  NOR4_X1 U569 ( .A1(n1274), .A2(n1275), .A3(n1276), .A4(n1277), .ZN(n1256) );
  NOR4_X1 U570 ( .A1(n1258), .A2(n1259), .A3(n1260), .A4(n1261), .ZN(n1257) );
  OAI221_X1 U571 ( .B1(n4725), .B2(n1287), .C1(n4723), .C2(n1288), .A(n1289), 
        .ZN(n1274) );
  NAND2_X1 U572 ( .A1(n1222), .A2(n1223), .ZN(N2507) );
  NOR4_X1 U573 ( .A1(n1240), .A2(n1241), .A3(n1242), .A4(n1243), .ZN(n1222) );
  NOR4_X1 U574 ( .A1(n1224), .A2(n1225), .A3(n1226), .A4(n1227), .ZN(n1223) );
  OAI221_X1 U575 ( .B1(n4726), .B2(n1253), .C1(n4723), .C2(n1254), .A(n1255), 
        .ZN(n1240) );
  NAND2_X1 U576 ( .A1(n1188), .A2(n1189), .ZN(N2509) );
  NOR4_X1 U577 ( .A1(n1206), .A2(n1207), .A3(n1208), .A4(n1209), .ZN(n1188) );
  NOR4_X1 U578 ( .A1(n1190), .A2(n1191), .A3(n1192), .A4(n1193), .ZN(n1189) );
  OAI221_X1 U579 ( .B1(n4726), .B2(n1219), .C1(n4723), .C2(n1220), .A(n1221), 
        .ZN(n1206) );
  NAND2_X1 U580 ( .A1(n1154), .A2(n1155), .ZN(N2511) );
  NOR4_X1 U581 ( .A1(n1172), .A2(n1173), .A3(n1174), .A4(n1175), .ZN(n1154) );
  NOR4_X1 U582 ( .A1(n1156), .A2(n1157), .A3(n1158), .A4(n1159), .ZN(n1155) );
  OAI221_X1 U583 ( .B1(n4726), .B2(n1185), .C1(n4723), .C2(n1186), .A(n1187), 
        .ZN(n1172) );
  NAND2_X1 U584 ( .A1(n1120), .A2(n1121), .ZN(N2513) );
  NOR4_X1 U585 ( .A1(n1138), .A2(n1139), .A3(n1140), .A4(n1141), .ZN(n1120) );
  NOR4_X1 U586 ( .A1(n1122), .A2(n1123), .A3(n1124), .A4(n1125), .ZN(n1121) );
  OAI221_X1 U587 ( .B1(n4726), .B2(n1151), .C1(n4723), .C2(n1152), .A(n1153), 
        .ZN(n1138) );
  NAND2_X1 U588 ( .A1(n1086), .A2(n1087), .ZN(N2515) );
  NOR4_X1 U589 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1086) );
  NOR4_X1 U590 ( .A1(n1088), .A2(n1089), .A3(n1090), .A4(n1091), .ZN(n1087) );
  OAI221_X1 U591 ( .B1(n4726), .B2(n1117), .C1(n4723), .C2(n1118), .A(n1119), 
        .ZN(n1104) );
  NAND2_X1 U592 ( .A1(n1052), .A2(n1053), .ZN(N2517) );
  NOR4_X1 U593 ( .A1(n1070), .A2(n1071), .A3(n1072), .A4(n1073), .ZN(n1052) );
  NOR4_X1 U594 ( .A1(n1054), .A2(n1055), .A3(n1056), .A4(n1057), .ZN(n1053) );
  OAI221_X1 U595 ( .B1(n4726), .B2(n1083), .C1(n4723), .C2(n1084), .A(n1085), 
        .ZN(n1070) );
  NAND2_X1 U596 ( .A1(n1018), .A2(n1019), .ZN(N2519) );
  NOR4_X1 U597 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1018) );
  NOR4_X1 U598 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1019) );
  OAI221_X1 U599 ( .B1(n4726), .B2(n1049), .C1(n4723), .C2(n1050), .A(n1051), 
        .ZN(n1036) );
  NAND2_X1 U600 ( .A1(n984), .A2(n985), .ZN(N2521) );
  NOR4_X1 U601 ( .A1(n1002), .A2(n1003), .A3(n1004), .A4(n1005), .ZN(n984) );
  NOR4_X1 U602 ( .A1(n986), .A2(n987), .A3(n988), .A4(n989), .ZN(n985) );
  OAI221_X1 U603 ( .B1(n4726), .B2(n1015), .C1(n4723), .C2(n1016), .A(n1017), 
        .ZN(n1002) );
  NAND2_X1 U604 ( .A1(n950), .A2(n951), .ZN(N2523) );
  NOR4_X1 U605 ( .A1(n968), .A2(n969), .A3(n970), .A4(n971), .ZN(n950) );
  NOR4_X1 U606 ( .A1(n952), .A2(n953), .A3(n954), .A4(n955), .ZN(n951) );
  OAI221_X1 U607 ( .B1(n4726), .B2(n981), .C1(n4723), .C2(n982), .A(n983), 
        .ZN(n968) );
  NAND2_X1 U608 ( .A1(n916), .A2(n917), .ZN(N2525) );
  NOR4_X1 U609 ( .A1(n934), .A2(n935), .A3(n936), .A4(n937), .ZN(n916) );
  NOR4_X1 U610 ( .A1(n918), .A2(n919), .A3(n920), .A4(n921), .ZN(n917) );
  OAI221_X1 U611 ( .B1(n4726), .B2(n947), .C1(n4723), .C2(n948), .A(n949), 
        .ZN(n934) );
  NAND2_X1 U612 ( .A1(n882), .A2(n883), .ZN(N2527) );
  NOR4_X1 U613 ( .A1(n900), .A2(n901), .A3(n902), .A4(n903), .ZN(n882) );
  NOR4_X1 U614 ( .A1(n884), .A2(n885), .A3(n886), .A4(n887), .ZN(n883) );
  OAI221_X1 U615 ( .B1(n4726), .B2(n913), .C1(n4724), .C2(n914), .A(n915), 
        .ZN(n900) );
  NAND2_X1 U616 ( .A1(n848), .A2(n849), .ZN(N2529) );
  NOR4_X1 U617 ( .A1(n866), .A2(n867), .A3(n868), .A4(n869), .ZN(n848) );
  NOR4_X1 U618 ( .A1(n850), .A2(n851), .A3(n852), .A4(n853), .ZN(n849) );
  OAI221_X1 U619 ( .B1(n4726), .B2(n879), .C1(n4724), .C2(n880), .A(n881), 
        .ZN(n866) );
  NAND2_X1 U620 ( .A1(n814), .A2(n815), .ZN(N2531) );
  NOR4_X1 U621 ( .A1(n832), .A2(n833), .A3(n834), .A4(n835), .ZN(n814) );
  NOR4_X1 U622 ( .A1(n816), .A2(n817), .A3(n818), .A4(n819), .ZN(n815) );
  OAI221_X1 U623 ( .B1(n4727), .B2(n845), .C1(n4724), .C2(n846), .A(n847), 
        .ZN(n832) );
  NAND2_X1 U624 ( .A1(n780), .A2(n781), .ZN(N2533) );
  NOR4_X1 U625 ( .A1(n798), .A2(n799), .A3(n800), .A4(n801), .ZN(n780) );
  NOR4_X1 U626 ( .A1(n782), .A2(n783), .A3(n784), .A4(n785), .ZN(n781) );
  OAI221_X1 U627 ( .B1(n4727), .B2(n811), .C1(n4724), .C2(n812), .A(n813), 
        .ZN(n798) );
  NAND2_X1 U628 ( .A1(n746), .A2(n747), .ZN(N2535) );
  NOR4_X1 U629 ( .A1(n764), .A2(n765), .A3(n766), .A4(n767), .ZN(n746) );
  NOR4_X1 U630 ( .A1(n748), .A2(n749), .A3(n750), .A4(n751), .ZN(n747) );
  OAI221_X1 U631 ( .B1(n4727), .B2(n777), .C1(n4724), .C2(n778), .A(n779), 
        .ZN(n764) );
  NAND2_X1 U632 ( .A1(n712), .A2(n713), .ZN(N2537) );
  NOR4_X1 U633 ( .A1(n730), .A2(n731), .A3(n732), .A4(n733), .ZN(n712) );
  NOR4_X1 U634 ( .A1(n714), .A2(n715), .A3(n716), .A4(n717), .ZN(n713) );
  OAI221_X1 U635 ( .B1(n4727), .B2(n743), .C1(n4724), .C2(n744), .A(n745), 
        .ZN(n730) );
  NAND2_X1 U636 ( .A1(n678), .A2(n679), .ZN(N2539) );
  NOR4_X1 U637 ( .A1(n696), .A2(n697), .A3(n698), .A4(n699), .ZN(n678) );
  NOR4_X1 U638 ( .A1(n680), .A2(n681), .A3(n682), .A4(n683), .ZN(n679) );
  OAI221_X1 U639 ( .B1(n4727), .B2(n709), .C1(n4724), .C2(n710), .A(n711), 
        .ZN(n696) );
  NAND2_X1 U640 ( .A1(n644), .A2(n645), .ZN(N2541) );
  NOR4_X1 U641 ( .A1(n662), .A2(n663), .A3(n664), .A4(n665), .ZN(n644) );
  NOR4_X1 U642 ( .A1(n646), .A2(n647), .A3(n648), .A4(n649), .ZN(n645) );
  OAI221_X1 U643 ( .B1(n4727), .B2(n675), .C1(n4724), .C2(n676), .A(n677), 
        .ZN(n662) );
  NAND2_X1 U644 ( .A1(n610), .A2(n611), .ZN(N2543) );
  NOR4_X1 U645 ( .A1(n628), .A2(n629), .A3(n630), .A4(n631), .ZN(n610) );
  NOR4_X1 U646 ( .A1(n612), .A2(n613), .A3(n614), .A4(n615), .ZN(n611) );
  OAI221_X1 U647 ( .B1(n4727), .B2(n641), .C1(n4724), .C2(n642), .A(n643), 
        .ZN(n628) );
  NAND2_X1 U648 ( .A1(n544), .A2(n545), .ZN(N2545) );
  NOR4_X1 U649 ( .A1(n578), .A2(n579), .A3(n580), .A4(n581), .ZN(n544) );
  NOR4_X1 U650 ( .A1(n546), .A2(n547), .A3(n548), .A4(n549), .ZN(n545) );
  OAI221_X1 U651 ( .B1(n4727), .B2(n604), .C1(n4724), .C2(n606), .A(n607), 
        .ZN(n578) );
  AND2_X1 U652 ( .A1(n2278), .A2(n2287), .ZN(n1699) );
  AND2_X1 U653 ( .A1(n2278), .A2(n2286), .ZN(n1700) );
  AND2_X1 U654 ( .A1(n2279), .A2(n2278), .ZN(n1689) );
  AND2_X1 U655 ( .A1(n2277), .A2(n2278), .ZN(n1690) );
  INV_X1 U656 ( .A(ADD_WR[4]), .ZN(n539) );
  INV_X1 U657 ( .A(ADD_WR[3]), .ZN(n537) );
  NOR3_X1 U658 ( .A1(n1648), .A2(ADD_RD2[4]), .A3(n1657), .ZN(n1665) );
  NOR3_X1 U659 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(n1657), .ZN(n1666) );
  NOR3_X1 U660 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(n1648), .ZN(n1673) );
  NOR3_X1 U661 ( .A1(ADD_RD2[3]), .A2(ADD_RD2[4]), .A3(ADD_RD2[0]), .ZN(n1674)
         );
  NOR3_X1 U662 ( .A1(n2284), .A2(ADD_RD1[4]), .A3(n2289), .ZN(n2295) );
  NOR3_X1 U663 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(n2289), .ZN(n2296) );
  NOR3_X1 U664 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(n2284), .ZN(n2299) );
  NOR3_X1 U665 ( .A1(ADD_RD1[3]), .A2(ADD_RD1[4]), .A3(ADD_RD1[0]), .ZN(n2300)
         );
  AND3_X1 U666 ( .A1(ADD_RD2[1]), .A2(n1675), .A3(ADD_RD2[2]), .ZN(n1642) );
  AND3_X1 U667 ( .A1(ADD_RD1[1]), .A2(n1675), .A3(ADD_RD1[2]), .ZN(n2280) );
  OAI221_X1 U668 ( .B1(n4811), .B2(n820), .C1(n4808), .C2(n821), .A(n822), 
        .ZN(n819) );
  AOI22_X1 U669 ( .A1(\REGISTERS[28][24] ), .A2(n4805), .B1(
        \REGISTERS[29][24] ), .B2(n4802), .ZN(n822) );
  OAI221_X1 U670 ( .B1(n4763), .B2(n836), .C1(n4760), .C2(n837), .A(n838), 
        .ZN(n835) );
  AOI22_X1 U671 ( .A1(\REGISTERS[12][24] ), .A2(n4757), .B1(
        \REGISTERS[13][24] ), .B2(n4754), .ZN(n838) );
  OAI221_X1 U672 ( .B1(n4811), .B2(n786), .C1(n4808), .C2(n787), .A(n788), 
        .ZN(n785) );
  AOI22_X1 U673 ( .A1(\REGISTERS[28][25] ), .A2(n4805), .B1(
        \REGISTERS[29][25] ), .B2(n4802), .ZN(n788) );
  OAI221_X1 U674 ( .B1(n4763), .B2(n802), .C1(n4760), .C2(n803), .A(n804), 
        .ZN(n801) );
  AOI22_X1 U675 ( .A1(\REGISTERS[12][25] ), .A2(n4757), .B1(
        \REGISTERS[13][25] ), .B2(n4754), .ZN(n804) );
  OAI221_X1 U676 ( .B1(n4811), .B2(n752), .C1(n4808), .C2(n753), .A(n754), 
        .ZN(n751) );
  AOI22_X1 U677 ( .A1(\REGISTERS[28][26] ), .A2(n4805), .B1(
        \REGISTERS[29][26] ), .B2(n4802), .ZN(n754) );
  OAI221_X1 U678 ( .B1(n4763), .B2(n768), .C1(n4760), .C2(n769), .A(n770), 
        .ZN(n767) );
  AOI22_X1 U679 ( .A1(\REGISTERS[12][26] ), .A2(n4757), .B1(
        \REGISTERS[13][26] ), .B2(n4754), .ZN(n770) );
  OAI221_X1 U680 ( .B1(n4811), .B2(n718), .C1(n4808), .C2(n719), .A(n720), 
        .ZN(n717) );
  AOI22_X1 U681 ( .A1(\REGISTERS[28][27] ), .A2(n4805), .B1(
        \REGISTERS[29][27] ), .B2(n4802), .ZN(n720) );
  OAI221_X1 U682 ( .B1(n4763), .B2(n734), .C1(n4760), .C2(n735), .A(n736), 
        .ZN(n733) );
  AOI22_X1 U683 ( .A1(\REGISTERS[12][27] ), .A2(n4757), .B1(
        \REGISTERS[13][27] ), .B2(n4754), .ZN(n736) );
  OAI221_X1 U684 ( .B1(n4811), .B2(n684), .C1(n4808), .C2(n685), .A(n686), 
        .ZN(n683) );
  AOI22_X1 U685 ( .A1(\REGISTERS[28][28] ), .A2(n4805), .B1(
        \REGISTERS[29][28] ), .B2(n4802), .ZN(n686) );
  OAI221_X1 U686 ( .B1(n4763), .B2(n700), .C1(n4760), .C2(n701), .A(n702), 
        .ZN(n699) );
  AOI22_X1 U687 ( .A1(\REGISTERS[12][28] ), .A2(n4757), .B1(
        \REGISTERS[13][28] ), .B2(n4754), .ZN(n702) );
  OAI221_X1 U688 ( .B1(n4811), .B2(n650), .C1(n4808), .C2(n651), .A(n652), 
        .ZN(n649) );
  AOI22_X1 U689 ( .A1(\REGISTERS[28][29] ), .A2(n4805), .B1(
        \REGISTERS[29][29] ), .B2(n4802), .ZN(n652) );
  OAI221_X1 U690 ( .B1(n4763), .B2(n666), .C1(n4760), .C2(n667), .A(n668), 
        .ZN(n665) );
  AOI22_X1 U691 ( .A1(\REGISTERS[12][29] ), .A2(n4757), .B1(
        \REGISTERS[13][29] ), .B2(n4754), .ZN(n668) );
  OAI221_X1 U692 ( .B1(n4811), .B2(n616), .C1(n4808), .C2(n617), .A(n618), 
        .ZN(n615) );
  AOI22_X1 U693 ( .A1(\REGISTERS[28][30] ), .A2(n4805), .B1(
        \REGISTERS[29][30] ), .B2(n4802), .ZN(n618) );
  OAI221_X1 U694 ( .B1(n4763), .B2(n632), .C1(n4760), .C2(n633), .A(n634), 
        .ZN(n631) );
  AOI22_X1 U695 ( .A1(\REGISTERS[12][30] ), .A2(n4757), .B1(
        \REGISTERS[13][30] ), .B2(n4754), .ZN(n634) );
  OAI221_X1 U696 ( .B1(n4811), .B2(n551), .C1(n4808), .C2(n553), .A(n554), 
        .ZN(n549) );
  AOI22_X1 U697 ( .A1(\REGISTERS[28][31] ), .A2(n4805), .B1(
        \REGISTERS[29][31] ), .B2(n4802), .ZN(n554) );
  OAI221_X1 U698 ( .B1(n4763), .B2(n583), .C1(n4760), .C2(n585), .A(n586), 
        .ZN(n581) );
  AOI22_X1 U699 ( .A1(\REGISTERS[12][31] ), .A2(n4757), .B1(
        \REGISTERS[13][31] ), .B2(n4754), .ZN(n586) );
  OAI221_X1 U700 ( .B1(n1636), .B2(n4713), .C1(n1637), .C2(n4710), .A(n2276), 
        .ZN(n2275) );
  AOI22_X1 U701 ( .A1(n4707), .A2(\REGISTERS[28][0] ), .B1(n4704), .B2(
        \REGISTERS[29][0] ), .ZN(n2276) );
  OAI221_X1 U702 ( .B1(n1662), .B2(n4665), .C1(n1663), .C2(n4662), .A(n2294), 
        .ZN(n2293) );
  AOI22_X1 U703 ( .A1(n4659), .A2(\REGISTERS[12][0] ), .B1(n4656), .B2(
        \REGISTERS[13][0] ), .ZN(n2294) );
  OAI221_X1 U704 ( .B1(n1602), .B2(n4713), .C1(n1603), .C2(n4710), .A(n2258), 
        .ZN(n2257) );
  AOI22_X1 U705 ( .A1(n4707), .A2(\REGISTERS[28][1] ), .B1(n4704), .B2(
        \REGISTERS[29][1] ), .ZN(n2258) );
  OAI221_X1 U706 ( .B1(n1618), .B2(n4665), .C1(n1619), .C2(n4662), .A(n2266), 
        .ZN(n2265) );
  AOI22_X1 U707 ( .A1(n4659), .A2(\REGISTERS[12][1] ), .B1(n4656), .B2(
        \REGISTERS[13][1] ), .ZN(n2266) );
  OAI221_X1 U708 ( .B1(n1568), .B2(n4713), .C1(n1569), .C2(n4710), .A(n2240), 
        .ZN(n2239) );
  AOI22_X1 U709 ( .A1(n4707), .A2(\REGISTERS[28][2] ), .B1(n4704), .B2(
        \REGISTERS[29][2] ), .ZN(n2240) );
  OAI221_X1 U710 ( .B1(n1584), .B2(n4665), .C1(n1585), .C2(n4662), .A(n2248), 
        .ZN(n2247) );
  AOI22_X1 U711 ( .A1(n4659), .A2(\REGISTERS[12][2] ), .B1(n4656), .B2(
        \REGISTERS[13][2] ), .ZN(n2248) );
  OAI221_X1 U712 ( .B1(n1534), .B2(n4713), .C1(n1535), .C2(n4710), .A(n2222), 
        .ZN(n2221) );
  AOI22_X1 U713 ( .A1(n4707), .A2(\REGISTERS[28][3] ), .B1(n4704), .B2(
        \REGISTERS[29][3] ), .ZN(n2222) );
  OAI221_X1 U714 ( .B1(n1550), .B2(n4665), .C1(n1551), .C2(n4662), .A(n2230), 
        .ZN(n2229) );
  AOI22_X1 U715 ( .A1(n4659), .A2(\REGISTERS[12][3] ), .B1(n4656), .B2(
        \REGISTERS[13][3] ), .ZN(n2230) );
  OAI221_X1 U716 ( .B1(n1500), .B2(n4713), .C1(n1501), .C2(n4710), .A(n2204), 
        .ZN(n2203) );
  AOI22_X1 U717 ( .A1(n4707), .A2(\REGISTERS[28][4] ), .B1(n4704), .B2(
        \REGISTERS[29][4] ), .ZN(n2204) );
  OAI221_X1 U718 ( .B1(n1516), .B2(n4665), .C1(n1517), .C2(n4662), .A(n2212), 
        .ZN(n2211) );
  AOI22_X1 U719 ( .A1(n4659), .A2(\REGISTERS[12][4] ), .B1(n4656), .B2(
        \REGISTERS[13][4] ), .ZN(n2212) );
  OAI221_X1 U720 ( .B1(n1466), .B2(n4713), .C1(n1467), .C2(n4710), .A(n2186), 
        .ZN(n2185) );
  AOI22_X1 U721 ( .A1(n4707), .A2(\REGISTERS[28][5] ), .B1(n4704), .B2(
        \REGISTERS[29][5] ), .ZN(n2186) );
  OAI221_X1 U722 ( .B1(n1482), .B2(n4665), .C1(n1483), .C2(n4662), .A(n2194), 
        .ZN(n2193) );
  AOI22_X1 U723 ( .A1(n4659), .A2(\REGISTERS[12][5] ), .B1(n4656), .B2(
        \REGISTERS[13][5] ), .ZN(n2194) );
  OAI221_X1 U724 ( .B1(n1432), .B2(n4713), .C1(n1433), .C2(n4710), .A(n2168), 
        .ZN(n2167) );
  AOI22_X1 U725 ( .A1(n4707), .A2(\REGISTERS[28][6] ), .B1(n4704), .B2(
        \REGISTERS[29][6] ), .ZN(n2168) );
  OAI221_X1 U726 ( .B1(n1448), .B2(n4665), .C1(n1449), .C2(n4662), .A(n2176), 
        .ZN(n2175) );
  AOI22_X1 U728 ( .A1(n4659), .A2(\REGISTERS[12][6] ), .B1(n4656), .B2(
        \REGISTERS[13][6] ), .ZN(n2176) );
  OAI221_X1 U729 ( .B1(n1398), .B2(n4713), .C1(n1399), .C2(n4710), .A(n2150), 
        .ZN(n2149) );
  AOI22_X1 U730 ( .A1(n4707), .A2(\REGISTERS[28][7] ), .B1(n4704), .B2(
        \REGISTERS[29][7] ), .ZN(n2150) );
  OAI221_X1 U731 ( .B1(n1414), .B2(n4665), .C1(n1415), .C2(n4662), .A(n2158), 
        .ZN(n2157) );
  AOI22_X1 U732 ( .A1(n4659), .A2(\REGISTERS[12][7] ), .B1(n4656), .B2(
        \REGISTERS[13][7] ), .ZN(n2158) );
  OAI221_X1 U733 ( .B1(n1364), .B2(n4713), .C1(n1365), .C2(n4710), .A(n2132), 
        .ZN(n2131) );
  AOI22_X1 U734 ( .A1(n4707), .A2(\REGISTERS[28][8] ), .B1(n4704), .B2(
        \REGISTERS[29][8] ), .ZN(n2132) );
  OAI221_X1 U735 ( .B1(n1380), .B2(n4665), .C1(n1381), .C2(n4662), .A(n2140), 
        .ZN(n2139) );
  AOI22_X1 U736 ( .A1(n4659), .A2(\REGISTERS[12][8] ), .B1(n4656), .B2(
        \REGISTERS[13][8] ), .ZN(n2140) );
  OAI221_X1 U737 ( .B1(n1330), .B2(n4713), .C1(n1331), .C2(n4710), .A(n2114), 
        .ZN(n2113) );
  AOI22_X1 U738 ( .A1(n4707), .A2(\REGISTERS[28][9] ), .B1(n4704), .B2(
        \REGISTERS[29][9] ), .ZN(n2114) );
  OAI221_X1 U739 ( .B1(n1346), .B2(n4665), .C1(n1347), .C2(n4662), .A(n2122), 
        .ZN(n2121) );
  AOI22_X1 U740 ( .A1(n4659), .A2(\REGISTERS[12][9] ), .B1(n4656), .B2(
        \REGISTERS[13][9] ), .ZN(n2122) );
  OAI221_X1 U741 ( .B1(n1296), .B2(n4713), .C1(n1297), .C2(n4710), .A(n2096), 
        .ZN(n2095) );
  AOI22_X1 U742 ( .A1(n4707), .A2(\REGISTERS[28][10] ), .B1(n4704), .B2(
        \REGISTERS[29][10] ), .ZN(n2096) );
  OAI221_X1 U743 ( .B1(n1312), .B2(n4665), .C1(n1313), .C2(n4662), .A(n2104), 
        .ZN(n2103) );
  AOI22_X1 U744 ( .A1(n4659), .A2(\REGISTERS[12][10] ), .B1(n4656), .B2(
        \REGISTERS[13][10] ), .ZN(n2104) );
  OAI221_X1 U745 ( .B1(n888), .B2(n4715), .C1(n889), .C2(n4712), .A(n1880), 
        .ZN(n1879) );
  AOI22_X1 U746 ( .A1(n4709), .A2(\REGISTERS[28][22] ), .B1(n4706), .B2(
        \REGISTERS[29][22] ), .ZN(n1880) );
  OAI221_X1 U747 ( .B1(n904), .B2(n4667), .C1(n905), .C2(n4664), .A(n1888), 
        .ZN(n1887) );
  AOI22_X1 U748 ( .A1(n4661), .A2(\REGISTERS[12][22] ), .B1(n4658), .B2(
        \REGISTERS[13][22] ), .ZN(n1888) );
  OAI221_X1 U749 ( .B1(n854), .B2(n4715), .C1(n855), .C2(n4712), .A(n1862), 
        .ZN(n1861) );
  AOI22_X1 U750 ( .A1(n4709), .A2(\REGISTERS[28][23] ), .B1(n4706), .B2(
        \REGISTERS[29][23] ), .ZN(n1862) );
  OAI221_X1 U751 ( .B1(n870), .B2(n4667), .C1(n871), .C2(n4664), .A(n1870), 
        .ZN(n1869) );
  AOI22_X1 U752 ( .A1(n4661), .A2(\REGISTERS[12][23] ), .B1(n4658), .B2(
        \REGISTERS[13][23] ), .ZN(n1870) );
  OAI221_X1 U753 ( .B1(n820), .B2(n4715), .C1(n821), .C2(n4712), .A(n1844), 
        .ZN(n1843) );
  AOI22_X1 U754 ( .A1(n4709), .A2(\REGISTERS[28][24] ), .B1(n4706), .B2(
        \REGISTERS[29][24] ), .ZN(n1844) );
  OAI221_X1 U755 ( .B1(n836), .B2(n4667), .C1(n837), .C2(n4664), .A(n1852), 
        .ZN(n1851) );
  AOI22_X1 U756 ( .A1(n4661), .A2(\REGISTERS[12][24] ), .B1(n4658), .B2(
        \REGISTERS[13][24] ), .ZN(n1852) );
  OAI221_X1 U757 ( .B1(n786), .B2(n4715), .C1(n787), .C2(n4712), .A(n1826), 
        .ZN(n1825) );
  AOI22_X1 U758 ( .A1(n4709), .A2(\REGISTERS[28][25] ), .B1(n4706), .B2(
        \REGISTERS[29][25] ), .ZN(n1826) );
  OAI221_X1 U759 ( .B1(n802), .B2(n4667), .C1(n803), .C2(n4664), .A(n1834), 
        .ZN(n1833) );
  AOI22_X1 U760 ( .A1(n4661), .A2(\REGISTERS[12][25] ), .B1(n4658), .B2(
        \REGISTERS[13][25] ), .ZN(n1834) );
  OAI221_X1 U761 ( .B1(n752), .B2(n4715), .C1(n753), .C2(n4712), .A(n1808), 
        .ZN(n1807) );
  AOI22_X1 U762 ( .A1(n4709), .A2(\REGISTERS[28][26] ), .B1(n4706), .B2(
        \REGISTERS[29][26] ), .ZN(n1808) );
  OAI221_X1 U763 ( .B1(n768), .B2(n4667), .C1(n769), .C2(n4664), .A(n1816), 
        .ZN(n1815) );
  AOI22_X1 U764 ( .A1(n4661), .A2(\REGISTERS[12][26] ), .B1(n4658), .B2(
        \REGISTERS[13][26] ), .ZN(n1816) );
  OAI221_X1 U765 ( .B1(n718), .B2(n4715), .C1(n719), .C2(n4712), .A(n1790), 
        .ZN(n1789) );
  AOI22_X1 U766 ( .A1(n4709), .A2(\REGISTERS[28][27] ), .B1(n4706), .B2(
        \REGISTERS[29][27] ), .ZN(n1790) );
  OAI221_X1 U767 ( .B1(n734), .B2(n4667), .C1(n735), .C2(n4664), .A(n1798), 
        .ZN(n1797) );
  AOI22_X1 U768 ( .A1(n4661), .A2(\REGISTERS[12][27] ), .B1(n4658), .B2(
        \REGISTERS[13][27] ), .ZN(n1798) );
  OAI221_X1 U769 ( .B1(n684), .B2(n4715), .C1(n685), .C2(n4712), .A(n1772), 
        .ZN(n1771) );
  AOI22_X1 U770 ( .A1(n4709), .A2(\REGISTERS[28][28] ), .B1(n4706), .B2(
        \REGISTERS[29][28] ), .ZN(n1772) );
  OAI221_X1 U771 ( .B1(n700), .B2(n4667), .C1(n701), .C2(n4664), .A(n1780), 
        .ZN(n1779) );
  AOI22_X1 U772 ( .A1(n4661), .A2(\REGISTERS[12][28] ), .B1(n4658), .B2(
        \REGISTERS[13][28] ), .ZN(n1780) );
  OAI221_X1 U773 ( .B1(n650), .B2(n4715), .C1(n651), .C2(n4712), .A(n1754), 
        .ZN(n1753) );
  AOI22_X1 U774 ( .A1(n4709), .A2(\REGISTERS[28][29] ), .B1(n4706), .B2(
        \REGISTERS[29][29] ), .ZN(n1754) );
  OAI221_X1 U775 ( .B1(n666), .B2(n4667), .C1(n667), .C2(n4664), .A(n1762), 
        .ZN(n1761) );
  AOI22_X1 U776 ( .A1(n4661), .A2(\REGISTERS[12][29] ), .B1(n4658), .B2(
        \REGISTERS[13][29] ), .ZN(n1762) );
  OAI221_X1 U777 ( .B1(n616), .B2(n4715), .C1(n617), .C2(n4712), .A(n1736), 
        .ZN(n1735) );
  AOI22_X1 U778 ( .A1(n4709), .A2(\REGISTERS[28][30] ), .B1(n4706), .B2(
        \REGISTERS[29][30] ), .ZN(n1736) );
  OAI221_X1 U779 ( .B1(n632), .B2(n4667), .C1(n633), .C2(n4664), .A(n1744), 
        .ZN(n1743) );
  AOI22_X1 U780 ( .A1(n4661), .A2(\REGISTERS[12][30] ), .B1(n4658), .B2(
        \REGISTERS[13][30] ), .ZN(n1744) );
  OAI221_X1 U781 ( .B1(n551), .B2(n4715), .C1(n553), .C2(n4712), .A(n1688), 
        .ZN(n1685) );
  AOI22_X1 U782 ( .A1(n4709), .A2(\REGISTERS[28][31] ), .B1(n4706), .B2(
        \REGISTERS[29][31] ), .ZN(n1688) );
  OAI221_X1 U783 ( .B1(n583), .B2(n4667), .C1(n585), .C2(n4664), .A(n1712), 
        .ZN(n1709) );
  AOI22_X1 U784 ( .A1(n4661), .A2(\REGISTERS[12][31] ), .B1(n4658), .B2(
        \REGISTERS[13][31] ), .ZN(n1712) );
  OAI221_X1 U785 ( .B1(n4799), .B2(n823), .C1(n4796), .C2(n824), .A(n825), 
        .ZN(n818) );
  AOI22_X1 U786 ( .A1(\REGISTERS[24][24] ), .A2(n4793), .B1(
        \REGISTERS[25][24] ), .B2(n4790), .ZN(n825) );
  OAI221_X1 U787 ( .B1(n4751), .B2(n839), .C1(n4748), .C2(n840), .A(n841), 
        .ZN(n834) );
  AOI22_X1 U788 ( .A1(\REGISTERS[8][24] ), .A2(n4745), .B1(\REGISTERS[9][24] ), 
        .B2(n4742), .ZN(n841) );
  OAI221_X1 U789 ( .B1(n4799), .B2(n789), .C1(n4796), .C2(n790), .A(n791), 
        .ZN(n784) );
  AOI22_X1 U790 ( .A1(\REGISTERS[24][25] ), .A2(n4793), .B1(
        \REGISTERS[25][25] ), .B2(n4790), .ZN(n791) );
  OAI221_X1 U791 ( .B1(n4751), .B2(n805), .C1(n4748), .C2(n806), .A(n807), 
        .ZN(n800) );
  AOI22_X1 U792 ( .A1(\REGISTERS[8][25] ), .A2(n4745), .B1(\REGISTERS[9][25] ), 
        .B2(n4742), .ZN(n807) );
  OAI221_X1 U793 ( .B1(n4799), .B2(n755), .C1(n4796), .C2(n756), .A(n757), 
        .ZN(n750) );
  AOI22_X1 U794 ( .A1(\REGISTERS[24][26] ), .A2(n4793), .B1(
        \REGISTERS[25][26] ), .B2(n4790), .ZN(n757) );
  OAI221_X1 U795 ( .B1(n4751), .B2(n771), .C1(n4748), .C2(n772), .A(n773), 
        .ZN(n766) );
  AOI22_X1 U796 ( .A1(\REGISTERS[8][26] ), .A2(n4745), .B1(\REGISTERS[9][26] ), 
        .B2(n4742), .ZN(n773) );
  OAI221_X1 U797 ( .B1(n4799), .B2(n721), .C1(n4796), .C2(n722), .A(n723), 
        .ZN(n716) );
  AOI22_X1 U798 ( .A1(\REGISTERS[24][27] ), .A2(n4793), .B1(
        \REGISTERS[25][27] ), .B2(n4790), .ZN(n723) );
  OAI221_X1 U799 ( .B1(n4751), .B2(n737), .C1(n4748), .C2(n738), .A(n739), 
        .ZN(n732) );
  AOI22_X1 U800 ( .A1(\REGISTERS[8][27] ), .A2(n4745), .B1(\REGISTERS[9][27] ), 
        .B2(n4742), .ZN(n739) );
  OAI221_X1 U801 ( .B1(n4799), .B2(n687), .C1(n4796), .C2(n688), .A(n689), 
        .ZN(n682) );
  AOI22_X1 U802 ( .A1(\REGISTERS[24][28] ), .A2(n4793), .B1(
        \REGISTERS[25][28] ), .B2(n4790), .ZN(n689) );
  OAI221_X1 U803 ( .B1(n4751), .B2(n703), .C1(n4748), .C2(n704), .A(n705), 
        .ZN(n698) );
  AOI22_X1 U804 ( .A1(\REGISTERS[8][28] ), .A2(n4745), .B1(\REGISTERS[9][28] ), 
        .B2(n4742), .ZN(n705) );
  OAI221_X1 U805 ( .B1(n4799), .B2(n653), .C1(n4796), .C2(n654), .A(n655), 
        .ZN(n648) );
  AOI22_X1 U806 ( .A1(\REGISTERS[24][29] ), .A2(n4793), .B1(
        \REGISTERS[25][29] ), .B2(n4790), .ZN(n655) );
  OAI221_X1 U807 ( .B1(n4751), .B2(n669), .C1(n4748), .C2(n670), .A(n671), 
        .ZN(n664) );
  AOI22_X1 U808 ( .A1(\REGISTERS[8][29] ), .A2(n4745), .B1(\REGISTERS[9][29] ), 
        .B2(n4742), .ZN(n671) );
  OAI221_X1 U809 ( .B1(n4799), .B2(n619), .C1(n4796), .C2(n620), .A(n621), 
        .ZN(n614) );
  AOI22_X1 U810 ( .A1(\REGISTERS[24][30] ), .A2(n4793), .B1(
        \REGISTERS[25][30] ), .B2(n4790), .ZN(n621) );
  OAI221_X1 U811 ( .B1(n4751), .B2(n635), .C1(n4748), .C2(n636), .A(n637), 
        .ZN(n630) );
  AOI22_X1 U812 ( .A1(\REGISTERS[8][30] ), .A2(n4745), .B1(\REGISTERS[9][30] ), 
        .B2(n4742), .ZN(n637) );
  OAI221_X1 U813 ( .B1(n4799), .B2(n558), .C1(n4796), .C2(n560), .A(n561), 
        .ZN(n548) );
  AOI22_X1 U814 ( .A1(\REGISTERS[24][31] ), .A2(n4793), .B1(
        \REGISTERS[25][31] ), .B2(n4790), .ZN(n561) );
  OAI221_X1 U815 ( .B1(n4751), .B2(n590), .C1(n4748), .C2(n592), .A(n593), 
        .ZN(n580) );
  AOI22_X1 U816 ( .A1(\REGISTERS[8][31] ), .A2(n4745), .B1(\REGISTERS[9][31] ), 
        .B2(n4742), .ZN(n593) );
  OAI221_X1 U817 ( .B1(n4809), .B2(n1636), .C1(n4806), .C2(n1637), .A(n1638), 
        .ZN(n1635) );
  AOI22_X1 U818 ( .A1(\REGISTERS[28][0] ), .A2(n4803), .B1(\REGISTERS[29][0] ), 
        .B2(n4800), .ZN(n1638) );
  OAI221_X1 U819 ( .B1(n4761), .B2(n1662), .C1(n4758), .C2(n1663), .A(n1664), 
        .ZN(n1661) );
  AOI22_X1 U820 ( .A1(\REGISTERS[12][0] ), .A2(n4755), .B1(\REGISTERS[13][0] ), 
        .B2(n4752), .ZN(n1664) );
  OAI221_X1 U821 ( .B1(n4809), .B2(n1602), .C1(n4806), .C2(n1603), .A(n1604), 
        .ZN(n1601) );
  AOI22_X1 U822 ( .A1(\REGISTERS[28][1] ), .A2(n4803), .B1(\REGISTERS[29][1] ), 
        .B2(n4800), .ZN(n1604) );
  OAI221_X1 U823 ( .B1(n4761), .B2(n1618), .C1(n4758), .C2(n1619), .A(n1620), 
        .ZN(n1617) );
  AOI22_X1 U824 ( .A1(\REGISTERS[12][1] ), .A2(n4755), .B1(\REGISTERS[13][1] ), 
        .B2(n4752), .ZN(n1620) );
  OAI221_X1 U825 ( .B1(n4809), .B2(n1568), .C1(n4806), .C2(n1569), .A(n1570), 
        .ZN(n1567) );
  AOI22_X1 U826 ( .A1(\REGISTERS[28][2] ), .A2(n4803), .B1(\REGISTERS[29][2] ), 
        .B2(n4800), .ZN(n1570) );
  OAI221_X1 U827 ( .B1(n4761), .B2(n1584), .C1(n4758), .C2(n1585), .A(n1586), 
        .ZN(n1583) );
  AOI22_X1 U828 ( .A1(\REGISTERS[12][2] ), .A2(n4755), .B1(\REGISTERS[13][2] ), 
        .B2(n4752), .ZN(n1586) );
  OAI221_X1 U829 ( .B1(n4809), .B2(n1534), .C1(n4806), .C2(n1535), .A(n1536), 
        .ZN(n1533) );
  AOI22_X1 U830 ( .A1(\REGISTERS[28][3] ), .A2(n4803), .B1(\REGISTERS[29][3] ), 
        .B2(n4800), .ZN(n1536) );
  OAI221_X1 U831 ( .B1(n4761), .B2(n1550), .C1(n4758), .C2(n1551), .A(n1552), 
        .ZN(n1549) );
  AOI22_X1 U832 ( .A1(\REGISTERS[12][3] ), .A2(n4755), .B1(\REGISTERS[13][3] ), 
        .B2(n4752), .ZN(n1552) );
  OAI221_X1 U833 ( .B1(n4809), .B2(n1500), .C1(n4806), .C2(n1501), .A(n1502), 
        .ZN(n1499) );
  AOI22_X1 U834 ( .A1(\REGISTERS[28][4] ), .A2(n4803), .B1(\REGISTERS[29][4] ), 
        .B2(n4800), .ZN(n1502) );
  OAI221_X1 U835 ( .B1(n4761), .B2(n1516), .C1(n4758), .C2(n1517), .A(n1518), 
        .ZN(n1515) );
  AOI22_X1 U836 ( .A1(\REGISTERS[12][4] ), .A2(n4755), .B1(\REGISTERS[13][4] ), 
        .B2(n4752), .ZN(n1518) );
  OAI221_X1 U837 ( .B1(n4809), .B2(n1466), .C1(n4806), .C2(n1467), .A(n1468), 
        .ZN(n1465) );
  AOI22_X1 U838 ( .A1(\REGISTERS[28][5] ), .A2(n4803), .B1(\REGISTERS[29][5] ), 
        .B2(n4800), .ZN(n1468) );
  OAI221_X1 U839 ( .B1(n4761), .B2(n1482), .C1(n4758), .C2(n1483), .A(n1484), 
        .ZN(n1481) );
  AOI22_X1 U840 ( .A1(\REGISTERS[12][5] ), .A2(n4755), .B1(\REGISTERS[13][5] ), 
        .B2(n4752), .ZN(n1484) );
  OAI221_X1 U841 ( .B1(n4809), .B2(n1432), .C1(n4806), .C2(n1433), .A(n1434), 
        .ZN(n1431) );
  AOI22_X1 U842 ( .A1(\REGISTERS[28][6] ), .A2(n4803), .B1(\REGISTERS[29][6] ), 
        .B2(n4800), .ZN(n1434) );
  OAI221_X1 U843 ( .B1(n4761), .B2(n1448), .C1(n4758), .C2(n1449), .A(n1450), 
        .ZN(n1447) );
  AOI22_X1 U844 ( .A1(\REGISTERS[12][6] ), .A2(n4755), .B1(\REGISTERS[13][6] ), 
        .B2(n4752), .ZN(n1450) );
  OAI221_X1 U845 ( .B1(n4809), .B2(n1398), .C1(n4806), .C2(n1399), .A(n1400), 
        .ZN(n1397) );
  AOI22_X1 U846 ( .A1(\REGISTERS[28][7] ), .A2(n4803), .B1(\REGISTERS[29][7] ), 
        .B2(n4800), .ZN(n1400) );
  OAI221_X1 U847 ( .B1(n4761), .B2(n1414), .C1(n4758), .C2(n1415), .A(n1416), 
        .ZN(n1413) );
  AOI22_X1 U848 ( .A1(\REGISTERS[12][7] ), .A2(n4755), .B1(\REGISTERS[13][7] ), 
        .B2(n4752), .ZN(n1416) );
  OAI221_X1 U849 ( .B1(n4809), .B2(n1364), .C1(n4806), .C2(n1365), .A(n1366), 
        .ZN(n1363) );
  AOI22_X1 U850 ( .A1(\REGISTERS[28][8] ), .A2(n4803), .B1(\REGISTERS[29][8] ), 
        .B2(n4800), .ZN(n1366) );
  OAI221_X1 U851 ( .B1(n4761), .B2(n1380), .C1(n4758), .C2(n1381), .A(n1382), 
        .ZN(n1379) );
  AOI22_X1 U852 ( .A1(\REGISTERS[12][8] ), .A2(n4755), .B1(\REGISTERS[13][8] ), 
        .B2(n4752), .ZN(n1382) );
  OAI221_X1 U853 ( .B1(n4809), .B2(n1330), .C1(n4806), .C2(n1331), .A(n1332), 
        .ZN(n1329) );
  AOI22_X1 U854 ( .A1(\REGISTERS[28][9] ), .A2(n4803), .B1(\REGISTERS[29][9] ), 
        .B2(n4800), .ZN(n1332) );
  OAI221_X1 U855 ( .B1(n4761), .B2(n1346), .C1(n4758), .C2(n1347), .A(n1348), 
        .ZN(n1345) );
  AOI22_X1 U856 ( .A1(\REGISTERS[12][9] ), .A2(n4755), .B1(\REGISTERS[13][9] ), 
        .B2(n4752), .ZN(n1348) );
  OAI221_X1 U857 ( .B1(n4809), .B2(n1296), .C1(n4806), .C2(n1297), .A(n1298), 
        .ZN(n1295) );
  AOI22_X1 U858 ( .A1(\REGISTERS[28][10] ), .A2(n4803), .B1(
        \REGISTERS[29][10] ), .B2(n4800), .ZN(n1298) );
  OAI221_X1 U859 ( .B1(n4761), .B2(n1312), .C1(n4758), .C2(n1313), .A(n1314), 
        .ZN(n1311) );
  AOI22_X1 U860 ( .A1(\REGISTERS[12][10] ), .A2(n4755), .B1(
        \REGISTERS[13][10] ), .B2(n4752), .ZN(n1314) );
  OAI221_X1 U861 ( .B1(n4809), .B2(n1262), .C1(n4807), .C2(n1263), .A(n1264), 
        .ZN(n1261) );
  AOI22_X1 U862 ( .A1(\REGISTERS[28][11] ), .A2(n4803), .B1(
        \REGISTERS[29][11] ), .B2(n4800), .ZN(n1264) );
  OAI221_X1 U863 ( .B1(n4761), .B2(n1278), .C1(n4759), .C2(n1279), .A(n1280), 
        .ZN(n1277) );
  AOI22_X1 U864 ( .A1(\REGISTERS[12][11] ), .A2(n4755), .B1(
        \REGISTERS[13][11] ), .B2(n4752), .ZN(n1280) );
  OAI221_X1 U865 ( .B1(n4810), .B2(n1228), .C1(n4807), .C2(n1229), .A(n1230), 
        .ZN(n1227) );
  AOI22_X1 U866 ( .A1(\REGISTERS[28][12] ), .A2(n4804), .B1(
        \REGISTERS[29][12] ), .B2(n4801), .ZN(n1230) );
  OAI221_X1 U867 ( .B1(n4762), .B2(n1244), .C1(n4759), .C2(n1245), .A(n1246), 
        .ZN(n1243) );
  AOI22_X1 U868 ( .A1(\REGISTERS[12][12] ), .A2(n4756), .B1(
        \REGISTERS[13][12] ), .B2(n4753), .ZN(n1246) );
  OAI221_X1 U869 ( .B1(n4810), .B2(n1194), .C1(n4807), .C2(n1195), .A(n1196), 
        .ZN(n1193) );
  AOI22_X1 U870 ( .A1(\REGISTERS[28][13] ), .A2(n4804), .B1(
        \REGISTERS[29][13] ), .B2(n4801), .ZN(n1196) );
  OAI221_X1 U871 ( .B1(n4762), .B2(n1210), .C1(n4759), .C2(n1211), .A(n1212), 
        .ZN(n1209) );
  AOI22_X1 U872 ( .A1(\REGISTERS[12][13] ), .A2(n4756), .B1(
        \REGISTERS[13][13] ), .B2(n4753), .ZN(n1212) );
  OAI221_X1 U873 ( .B1(n4810), .B2(n1160), .C1(n4807), .C2(n1161), .A(n1162), 
        .ZN(n1159) );
  AOI22_X1 U874 ( .A1(\REGISTERS[28][14] ), .A2(n4804), .B1(
        \REGISTERS[29][14] ), .B2(n4801), .ZN(n1162) );
  OAI221_X1 U875 ( .B1(n4762), .B2(n1176), .C1(n4759), .C2(n1177), .A(n1178), 
        .ZN(n1175) );
  AOI22_X1 U876 ( .A1(\REGISTERS[12][14] ), .A2(n4756), .B1(
        \REGISTERS[13][14] ), .B2(n4753), .ZN(n1178) );
  OAI221_X1 U877 ( .B1(n4810), .B2(n1126), .C1(n4807), .C2(n1127), .A(n1128), 
        .ZN(n1125) );
  AOI22_X1 U878 ( .A1(\REGISTERS[28][15] ), .A2(n4804), .B1(
        \REGISTERS[29][15] ), .B2(n4801), .ZN(n1128) );
  OAI221_X1 U879 ( .B1(n4762), .B2(n1142), .C1(n4759), .C2(n1143), .A(n1144), 
        .ZN(n1141) );
  AOI22_X1 U880 ( .A1(\REGISTERS[12][15] ), .A2(n4756), .B1(
        \REGISTERS[13][15] ), .B2(n4753), .ZN(n1144) );
  OAI221_X1 U881 ( .B1(n4810), .B2(n1092), .C1(n4807), .C2(n1093), .A(n1094), 
        .ZN(n1091) );
  AOI22_X1 U882 ( .A1(\REGISTERS[28][16] ), .A2(n4804), .B1(
        \REGISTERS[29][16] ), .B2(n4801), .ZN(n1094) );
  OAI221_X1 U883 ( .B1(n4762), .B2(n1108), .C1(n4759), .C2(n1109), .A(n1110), 
        .ZN(n1107) );
  AOI22_X1 U884 ( .A1(\REGISTERS[12][16] ), .A2(n4756), .B1(
        \REGISTERS[13][16] ), .B2(n4753), .ZN(n1110) );
  OAI221_X1 U885 ( .B1(n4810), .B2(n1058), .C1(n4807), .C2(n1059), .A(n1060), 
        .ZN(n1057) );
  AOI22_X1 U886 ( .A1(\REGISTERS[28][17] ), .A2(n4804), .B1(
        \REGISTERS[29][17] ), .B2(n4801), .ZN(n1060) );
  OAI221_X1 U887 ( .B1(n4762), .B2(n1074), .C1(n4759), .C2(n1075), .A(n1076), 
        .ZN(n1073) );
  AOI22_X1 U888 ( .A1(\REGISTERS[12][17] ), .A2(n4756), .B1(
        \REGISTERS[13][17] ), .B2(n4753), .ZN(n1076) );
  OAI221_X1 U889 ( .B1(n4810), .B2(n1024), .C1(n4807), .C2(n1025), .A(n1026), 
        .ZN(n1023) );
  AOI22_X1 U890 ( .A1(\REGISTERS[28][18] ), .A2(n4804), .B1(
        \REGISTERS[29][18] ), .B2(n4801), .ZN(n1026) );
  OAI221_X1 U891 ( .B1(n4762), .B2(n1040), .C1(n4759), .C2(n1041), .A(n1042), 
        .ZN(n1039) );
  AOI22_X1 U892 ( .A1(\REGISTERS[12][18] ), .A2(n4756), .B1(
        \REGISTERS[13][18] ), .B2(n4753), .ZN(n1042) );
  OAI221_X1 U893 ( .B1(n4810), .B2(n990), .C1(n4807), .C2(n991), .A(n992), 
        .ZN(n989) );
  AOI22_X1 U894 ( .A1(\REGISTERS[28][19] ), .A2(n4804), .B1(
        \REGISTERS[29][19] ), .B2(n4801), .ZN(n992) );
  OAI221_X1 U895 ( .B1(n4762), .B2(n1006), .C1(n4759), .C2(n1007), .A(n1008), 
        .ZN(n1005) );
  AOI22_X1 U896 ( .A1(\REGISTERS[12][19] ), .A2(n4756), .B1(
        \REGISTERS[13][19] ), .B2(n4753), .ZN(n1008) );
  OAI221_X1 U897 ( .B1(n4810), .B2(n956), .C1(n4807), .C2(n957), .A(n958), 
        .ZN(n955) );
  AOI22_X1 U898 ( .A1(\REGISTERS[28][20] ), .A2(n4804), .B1(
        \REGISTERS[29][20] ), .B2(n4801), .ZN(n958) );
  OAI221_X1 U899 ( .B1(n4762), .B2(n972), .C1(n4759), .C2(n973), .A(n974), 
        .ZN(n971) );
  AOI22_X1 U900 ( .A1(\REGISTERS[12][20] ), .A2(n4756), .B1(
        \REGISTERS[13][20] ), .B2(n4753), .ZN(n974) );
  OAI221_X1 U901 ( .B1(n4810), .B2(n922), .C1(n4807), .C2(n923), .A(n924), 
        .ZN(n921) );
  AOI22_X1 U902 ( .A1(\REGISTERS[28][21] ), .A2(n4804), .B1(
        \REGISTERS[29][21] ), .B2(n4801), .ZN(n924) );
  OAI221_X1 U903 ( .B1(n4762), .B2(n938), .C1(n4759), .C2(n939), .A(n940), 
        .ZN(n937) );
  AOI22_X1 U904 ( .A1(\REGISTERS[12][21] ), .A2(n4756), .B1(
        \REGISTERS[13][21] ), .B2(n4753), .ZN(n940) );
  OAI221_X1 U905 ( .B1(n4810), .B2(n888), .C1(n4808), .C2(n889), .A(n890), 
        .ZN(n887) );
  AOI22_X1 U906 ( .A1(\REGISTERS[28][22] ), .A2(n4804), .B1(
        \REGISTERS[29][22] ), .B2(n4801), .ZN(n890) );
  OAI221_X1 U907 ( .B1(n4762), .B2(n904), .C1(n4760), .C2(n905), .A(n906), 
        .ZN(n903) );
  AOI22_X1 U908 ( .A1(\REGISTERS[12][22] ), .A2(n4756), .B1(
        \REGISTERS[13][22] ), .B2(n4753), .ZN(n906) );
  OAI221_X1 U909 ( .B1(n4810), .B2(n854), .C1(n4808), .C2(n855), .A(n856), 
        .ZN(n853) );
  AOI22_X1 U910 ( .A1(\REGISTERS[28][23] ), .A2(n4804), .B1(
        \REGISTERS[29][23] ), .B2(n4801), .ZN(n856) );
  OAI221_X1 U911 ( .B1(n4762), .B2(n870), .C1(n4760), .C2(n871), .A(n872), 
        .ZN(n869) );
  AOI22_X1 U912 ( .A1(\REGISTERS[12][23] ), .A2(n4756), .B1(
        \REGISTERS[13][23] ), .B2(n4753), .ZN(n872) );
  OAI221_X1 U913 ( .B1(n1262), .B2(n4714), .C1(n1263), .C2(n4711), .A(n2078), 
        .ZN(n2077) );
  AOI22_X1 U914 ( .A1(n4708), .A2(\REGISTERS[28][11] ), .B1(n4705), .B2(
        \REGISTERS[29][11] ), .ZN(n2078) );
  OAI221_X1 U915 ( .B1(n1278), .B2(n4666), .C1(n1279), .C2(n4663), .A(n2086), 
        .ZN(n2085) );
  AOI22_X1 U916 ( .A1(n4660), .A2(\REGISTERS[12][11] ), .B1(n4657), .B2(
        \REGISTERS[13][11] ), .ZN(n2086) );
  OAI221_X1 U917 ( .B1(n1228), .B2(n4714), .C1(n1229), .C2(n4711), .A(n2060), 
        .ZN(n2059) );
  AOI22_X1 U918 ( .A1(n4708), .A2(\REGISTERS[28][12] ), .B1(n4705), .B2(
        \REGISTERS[29][12] ), .ZN(n2060) );
  OAI221_X1 U919 ( .B1(n1244), .B2(n4666), .C1(n1245), .C2(n4663), .A(n2068), 
        .ZN(n2067) );
  AOI22_X1 U920 ( .A1(n4660), .A2(\REGISTERS[12][12] ), .B1(n4657), .B2(
        \REGISTERS[13][12] ), .ZN(n2068) );
  OAI221_X1 U921 ( .B1(n1194), .B2(n4714), .C1(n1195), .C2(n4711), .A(n2042), 
        .ZN(n2041) );
  AOI22_X1 U922 ( .A1(n4708), .A2(\REGISTERS[28][13] ), .B1(n4705), .B2(
        \REGISTERS[29][13] ), .ZN(n2042) );
  OAI221_X1 U923 ( .B1(n1210), .B2(n4666), .C1(n1211), .C2(n4663), .A(n2050), 
        .ZN(n2049) );
  AOI22_X1 U924 ( .A1(n4660), .A2(\REGISTERS[12][13] ), .B1(n4657), .B2(
        \REGISTERS[13][13] ), .ZN(n2050) );
  OAI221_X1 U925 ( .B1(n1160), .B2(n4714), .C1(n1161), .C2(n4711), .A(n2024), 
        .ZN(n2023) );
  AOI22_X1 U926 ( .A1(n4708), .A2(\REGISTERS[28][14] ), .B1(n4705), .B2(
        \REGISTERS[29][14] ), .ZN(n2024) );
  OAI221_X1 U927 ( .B1(n1176), .B2(n4666), .C1(n1177), .C2(n4663), .A(n2032), 
        .ZN(n2031) );
  AOI22_X1 U928 ( .A1(n4660), .A2(\REGISTERS[12][14] ), .B1(n4657), .B2(
        \REGISTERS[13][14] ), .ZN(n2032) );
  OAI221_X1 U929 ( .B1(n1126), .B2(n4714), .C1(n1127), .C2(n4711), .A(n2006), 
        .ZN(n2005) );
  AOI22_X1 U930 ( .A1(n4708), .A2(\REGISTERS[28][15] ), .B1(n4705), .B2(
        \REGISTERS[29][15] ), .ZN(n2006) );
  OAI221_X1 U931 ( .B1(n1142), .B2(n4666), .C1(n1143), .C2(n4663), .A(n2014), 
        .ZN(n2013) );
  AOI22_X1 U932 ( .A1(n4660), .A2(\REGISTERS[12][15] ), .B1(n4657), .B2(
        \REGISTERS[13][15] ), .ZN(n2014) );
  OAI221_X1 U933 ( .B1(n1092), .B2(n4714), .C1(n1093), .C2(n4711), .A(n1988), 
        .ZN(n1987) );
  AOI22_X1 U934 ( .A1(n4708), .A2(\REGISTERS[28][16] ), .B1(n4705), .B2(
        \REGISTERS[29][16] ), .ZN(n1988) );
  OAI221_X1 U935 ( .B1(n1108), .B2(n4666), .C1(n1109), .C2(n4663), .A(n1996), 
        .ZN(n1995) );
  AOI22_X1 U936 ( .A1(n4660), .A2(\REGISTERS[12][16] ), .B1(n4657), .B2(
        \REGISTERS[13][16] ), .ZN(n1996) );
  OAI221_X1 U937 ( .B1(n1058), .B2(n4714), .C1(n1059), .C2(n4711), .A(n1970), 
        .ZN(n1969) );
  AOI22_X1 U938 ( .A1(n4708), .A2(\REGISTERS[28][17] ), .B1(n4705), .B2(
        \REGISTERS[29][17] ), .ZN(n1970) );
  OAI221_X1 U939 ( .B1(n1074), .B2(n4666), .C1(n1075), .C2(n4663), .A(n1978), 
        .ZN(n1977) );
  AOI22_X1 U940 ( .A1(n4660), .A2(\REGISTERS[12][17] ), .B1(n4657), .B2(
        \REGISTERS[13][17] ), .ZN(n1978) );
  OAI221_X1 U941 ( .B1(n1024), .B2(n4714), .C1(n1025), .C2(n4711), .A(n1952), 
        .ZN(n1951) );
  AOI22_X1 U942 ( .A1(n4708), .A2(\REGISTERS[28][18] ), .B1(n4705), .B2(
        \REGISTERS[29][18] ), .ZN(n1952) );
  OAI221_X1 U943 ( .B1(n1040), .B2(n4666), .C1(n1041), .C2(n4663), .A(n1960), 
        .ZN(n1959) );
  AOI22_X1 U944 ( .A1(n4660), .A2(\REGISTERS[12][18] ), .B1(n4657), .B2(
        \REGISTERS[13][18] ), .ZN(n1960) );
  OAI221_X1 U945 ( .B1(n990), .B2(n4714), .C1(n991), .C2(n4711), .A(n1934), 
        .ZN(n1933) );
  AOI22_X1 U946 ( .A1(n4708), .A2(\REGISTERS[28][19] ), .B1(n4705), .B2(
        \REGISTERS[29][19] ), .ZN(n1934) );
  OAI221_X1 U947 ( .B1(n1006), .B2(n4666), .C1(n1007), .C2(n4663), .A(n1942), 
        .ZN(n1941) );
  AOI22_X1 U948 ( .A1(n4660), .A2(\REGISTERS[12][19] ), .B1(n4657), .B2(
        \REGISTERS[13][19] ), .ZN(n1942) );
  OAI221_X1 U949 ( .B1(n956), .B2(n4714), .C1(n957), .C2(n4711), .A(n1916), 
        .ZN(n1915) );
  AOI22_X1 U950 ( .A1(n4708), .A2(\REGISTERS[28][20] ), .B1(n4705), .B2(
        \REGISTERS[29][20] ), .ZN(n1916) );
  OAI221_X1 U951 ( .B1(n972), .B2(n4666), .C1(n973), .C2(n4663), .A(n1924), 
        .ZN(n1923) );
  AOI22_X1 U952 ( .A1(n4660), .A2(\REGISTERS[12][20] ), .B1(n4657), .B2(
        \REGISTERS[13][20] ), .ZN(n1924) );
  OAI221_X1 U953 ( .B1(n922), .B2(n4714), .C1(n923), .C2(n4711), .A(n1898), 
        .ZN(n1897) );
  AOI22_X1 U954 ( .A1(n4708), .A2(\REGISTERS[28][21] ), .B1(n4705), .B2(
        \REGISTERS[29][21] ), .ZN(n1898) );
  OAI221_X1 U955 ( .B1(n938), .B2(n4666), .C1(n939), .C2(n4663), .A(n1906), 
        .ZN(n1905) );
  AOI22_X1 U956 ( .A1(n4660), .A2(\REGISTERS[12][21] ), .B1(n4657), .B2(
        \REGISTERS[13][21] ), .ZN(n1906) );
  OAI221_X1 U957 ( .B1(n1643), .B2(n4701), .C1(n1644), .C2(n4698), .A(n2281), 
        .ZN(n2274) );
  AOI22_X1 U958 ( .A1(n4695), .A2(\REGISTERS[24][0] ), .B1(n4692), .B2(
        \REGISTERS[25][0] ), .ZN(n2281) );
  OAI221_X1 U959 ( .B1(n1667), .B2(n4653), .C1(n1668), .C2(n4650), .A(n2297), 
        .ZN(n2292) );
  AOI22_X1 U960 ( .A1(n4647), .A2(\REGISTERS[8][0] ), .B1(n4644), .B2(
        \REGISTERS[9][0] ), .ZN(n2297) );
  OAI221_X1 U961 ( .B1(n1605), .B2(n4701), .C1(n1606), .C2(n4698), .A(n2259), 
        .ZN(n2256) );
  AOI22_X1 U962 ( .A1(n4695), .A2(\REGISTERS[24][1] ), .B1(n4692), .B2(
        \REGISTERS[25][1] ), .ZN(n2259) );
  OAI221_X1 U963 ( .B1(n1621), .B2(n4653), .C1(n1622), .C2(n4650), .A(n2267), 
        .ZN(n2264) );
  AOI22_X1 U964 ( .A1(n4647), .A2(\REGISTERS[8][1] ), .B1(n4644), .B2(
        \REGISTERS[9][1] ), .ZN(n2267) );
  OAI221_X1 U965 ( .B1(n1571), .B2(n4701), .C1(n1572), .C2(n4698), .A(n2241), 
        .ZN(n2238) );
  AOI22_X1 U966 ( .A1(n4695), .A2(\REGISTERS[24][2] ), .B1(n4692), .B2(
        \REGISTERS[25][2] ), .ZN(n2241) );
  OAI221_X1 U967 ( .B1(n1587), .B2(n4653), .C1(n1588), .C2(n4650), .A(n2249), 
        .ZN(n2246) );
  AOI22_X1 U968 ( .A1(n4647), .A2(\REGISTERS[8][2] ), .B1(n4644), .B2(
        \REGISTERS[9][2] ), .ZN(n2249) );
  OAI221_X1 U969 ( .B1(n1537), .B2(n4701), .C1(n1538), .C2(n4698), .A(n2223), 
        .ZN(n2220) );
  AOI22_X1 U970 ( .A1(n4695), .A2(\REGISTERS[24][3] ), .B1(n4692), .B2(
        \REGISTERS[25][3] ), .ZN(n2223) );
  OAI221_X1 U971 ( .B1(n1553), .B2(n4653), .C1(n1554), .C2(n4650), .A(n2231), 
        .ZN(n2228) );
  AOI22_X1 U972 ( .A1(n4647), .A2(\REGISTERS[8][3] ), .B1(n4644), .B2(
        \REGISTERS[9][3] ), .ZN(n2231) );
  OAI221_X1 U973 ( .B1(n1503), .B2(n4701), .C1(n1504), .C2(n4698), .A(n2205), 
        .ZN(n2202) );
  AOI22_X1 U974 ( .A1(n4695), .A2(\REGISTERS[24][4] ), .B1(n4692), .B2(
        \REGISTERS[25][4] ), .ZN(n2205) );
  OAI221_X1 U975 ( .B1(n1519), .B2(n4653), .C1(n1520), .C2(n4650), .A(n2213), 
        .ZN(n2210) );
  AOI22_X1 U976 ( .A1(n4647), .A2(\REGISTERS[8][4] ), .B1(n4644), .B2(
        \REGISTERS[9][4] ), .ZN(n2213) );
  OAI221_X1 U977 ( .B1(n1469), .B2(n4701), .C1(n1470), .C2(n4698), .A(n2187), 
        .ZN(n2184) );
  AOI22_X1 U978 ( .A1(n4695), .A2(\REGISTERS[24][5] ), .B1(n4692), .B2(
        \REGISTERS[25][5] ), .ZN(n2187) );
  OAI221_X1 U979 ( .B1(n1485), .B2(n4653), .C1(n1486), .C2(n4650), .A(n2195), 
        .ZN(n2192) );
  AOI22_X1 U980 ( .A1(n4647), .A2(\REGISTERS[8][5] ), .B1(n4644), .B2(
        \REGISTERS[9][5] ), .ZN(n2195) );
  OAI221_X1 U981 ( .B1(n1435), .B2(n4701), .C1(n1436), .C2(n4698), .A(n2169), 
        .ZN(n2166) );
  AOI22_X1 U982 ( .A1(n4695), .A2(\REGISTERS[24][6] ), .B1(n4692), .B2(
        \REGISTERS[25][6] ), .ZN(n2169) );
  OAI221_X1 U983 ( .B1(n1451), .B2(n4653), .C1(n1452), .C2(n4650), .A(n2177), 
        .ZN(n2174) );
  AOI22_X1 U984 ( .A1(n4647), .A2(\REGISTERS[8][6] ), .B1(n4644), .B2(
        \REGISTERS[9][6] ), .ZN(n2177) );
  OAI221_X1 U985 ( .B1(n1401), .B2(n4701), .C1(n1402), .C2(n4698), .A(n2151), 
        .ZN(n2148) );
  AOI22_X1 U986 ( .A1(n4695), .A2(\REGISTERS[24][7] ), .B1(n4692), .B2(
        \REGISTERS[25][7] ), .ZN(n2151) );
  OAI221_X1 U987 ( .B1(n1417), .B2(n4653), .C1(n1418), .C2(n4650), .A(n2159), 
        .ZN(n2156) );
  AOI22_X1 U988 ( .A1(n4647), .A2(\REGISTERS[8][7] ), .B1(n4644), .B2(
        \REGISTERS[9][7] ), .ZN(n2159) );
  OAI221_X1 U989 ( .B1(n1367), .B2(n4701), .C1(n1368), .C2(n4698), .A(n2133), 
        .ZN(n2130) );
  AOI22_X1 U990 ( .A1(n4695), .A2(\REGISTERS[24][8] ), .B1(n4692), .B2(
        \REGISTERS[25][8] ), .ZN(n2133) );
  OAI221_X1 U991 ( .B1(n1383), .B2(n4653), .C1(n1384), .C2(n4650), .A(n2141), 
        .ZN(n2138) );
  AOI22_X1 U992 ( .A1(n4647), .A2(\REGISTERS[8][8] ), .B1(n4644), .B2(
        \REGISTERS[9][8] ), .ZN(n2141) );
  OAI221_X1 U993 ( .B1(n1333), .B2(n4701), .C1(n1334), .C2(n4698), .A(n2115), 
        .ZN(n2112) );
  AOI22_X1 U994 ( .A1(n4695), .A2(\REGISTERS[24][9] ), .B1(n4692), .B2(
        \REGISTERS[25][9] ), .ZN(n2115) );
  OAI221_X1 U995 ( .B1(n1349), .B2(n4653), .C1(n1350), .C2(n4650), .A(n2123), 
        .ZN(n2120) );
  AOI22_X1 U996 ( .A1(n4647), .A2(\REGISTERS[8][9] ), .B1(n4644), .B2(
        \REGISTERS[9][9] ), .ZN(n2123) );
  OAI221_X1 U997 ( .B1(n1299), .B2(n4701), .C1(n1300), .C2(n4698), .A(n2097), 
        .ZN(n2094) );
  AOI22_X1 U998 ( .A1(n4695), .A2(\REGISTERS[24][10] ), .B1(n4692), .B2(
        \REGISTERS[25][10] ), .ZN(n2097) );
  OAI221_X1 U999 ( .B1(n1315), .B2(n4653), .C1(n1316), .C2(n4650), .A(n2105), 
        .ZN(n2102) );
  AOI22_X1 U1000 ( .A1(n4647), .A2(\REGISTERS[8][10] ), .B1(n4644), .B2(
        \REGISTERS[9][10] ), .ZN(n2105) );
  OAI221_X1 U1001 ( .B1(n891), .B2(n4703), .C1(n892), .C2(n4700), .A(n1881), 
        .ZN(n1878) );
  AOI22_X1 U1002 ( .A1(n4697), .A2(\REGISTERS[24][22] ), .B1(n4694), .B2(
        \REGISTERS[25][22] ), .ZN(n1881) );
  OAI221_X1 U1003 ( .B1(n907), .B2(n4655), .C1(n908), .C2(n4652), .A(n1889), 
        .ZN(n1886) );
  AOI22_X1 U1004 ( .A1(n4649), .A2(\REGISTERS[8][22] ), .B1(n4646), .B2(
        \REGISTERS[9][22] ), .ZN(n1889) );
  OAI221_X1 U1005 ( .B1(n857), .B2(n4703), .C1(n858), .C2(n4700), .A(n1863), 
        .ZN(n1860) );
  AOI22_X1 U1006 ( .A1(n4697), .A2(\REGISTERS[24][23] ), .B1(n4694), .B2(
        \REGISTERS[25][23] ), .ZN(n1863) );
  OAI221_X1 U1007 ( .B1(n873), .B2(n4655), .C1(n874), .C2(n4652), .A(n1871), 
        .ZN(n1868) );
  AOI22_X1 U1008 ( .A1(n4649), .A2(\REGISTERS[8][23] ), .B1(n4646), .B2(
        \REGISTERS[9][23] ), .ZN(n1871) );
  OAI221_X1 U1009 ( .B1(n823), .B2(n4703), .C1(n824), .C2(n4700), .A(n1845), 
        .ZN(n1842) );
  AOI22_X1 U1010 ( .A1(n4697), .A2(\REGISTERS[24][24] ), .B1(n4694), .B2(
        \REGISTERS[25][24] ), .ZN(n1845) );
  OAI221_X1 U1011 ( .B1(n839), .B2(n4655), .C1(n840), .C2(n4652), .A(n1853), 
        .ZN(n1850) );
  AOI22_X1 U1012 ( .A1(n4649), .A2(\REGISTERS[8][24] ), .B1(n4646), .B2(
        \REGISTERS[9][24] ), .ZN(n1853) );
  OAI221_X1 U1013 ( .B1(n789), .B2(n4703), .C1(n790), .C2(n4700), .A(n1827), 
        .ZN(n1824) );
  AOI22_X1 U1014 ( .A1(n4697), .A2(\REGISTERS[24][25] ), .B1(n4694), .B2(
        \REGISTERS[25][25] ), .ZN(n1827) );
  OAI221_X1 U1015 ( .B1(n805), .B2(n4655), .C1(n806), .C2(n4652), .A(n1835), 
        .ZN(n1832) );
  AOI22_X1 U1016 ( .A1(n4649), .A2(\REGISTERS[8][25] ), .B1(n4646), .B2(
        \REGISTERS[9][25] ), .ZN(n1835) );
  OAI221_X1 U1017 ( .B1(n755), .B2(n4703), .C1(n756), .C2(n4700), .A(n1809), 
        .ZN(n1806) );
  AOI22_X1 U1018 ( .A1(n4697), .A2(\REGISTERS[24][26] ), .B1(n4694), .B2(
        \REGISTERS[25][26] ), .ZN(n1809) );
  OAI221_X1 U1019 ( .B1(n771), .B2(n4655), .C1(n772), .C2(n4652), .A(n1817), 
        .ZN(n1814) );
  AOI22_X1 U1020 ( .A1(n4649), .A2(\REGISTERS[8][26] ), .B1(n4646), .B2(
        \REGISTERS[9][26] ), .ZN(n1817) );
  OAI221_X1 U1021 ( .B1(n721), .B2(n4703), .C1(n722), .C2(n4700), .A(n1791), 
        .ZN(n1788) );
  AOI22_X1 U1022 ( .A1(n4697), .A2(\REGISTERS[24][27] ), .B1(n4694), .B2(
        \REGISTERS[25][27] ), .ZN(n1791) );
  OAI221_X1 U1023 ( .B1(n737), .B2(n4655), .C1(n738), .C2(n4652), .A(n1799), 
        .ZN(n1796) );
  AOI22_X1 U1024 ( .A1(n4649), .A2(\REGISTERS[8][27] ), .B1(n4646), .B2(
        \REGISTERS[9][27] ), .ZN(n1799) );
  OAI221_X1 U1025 ( .B1(n687), .B2(n4703), .C1(n688), .C2(n4700), .A(n1773), 
        .ZN(n1770) );
  AOI22_X1 U1026 ( .A1(n4697), .A2(\REGISTERS[24][28] ), .B1(n4694), .B2(
        \REGISTERS[25][28] ), .ZN(n1773) );
  OAI221_X1 U1027 ( .B1(n703), .B2(n4655), .C1(n704), .C2(n4652), .A(n1781), 
        .ZN(n1778) );
  AOI22_X1 U1028 ( .A1(n4649), .A2(\REGISTERS[8][28] ), .B1(n4646), .B2(
        \REGISTERS[9][28] ), .ZN(n1781) );
  OAI221_X1 U1029 ( .B1(n653), .B2(n4703), .C1(n654), .C2(n4700), .A(n1755), 
        .ZN(n1752) );
  AOI22_X1 U1030 ( .A1(n4697), .A2(\REGISTERS[24][29] ), .B1(n4694), .B2(
        \REGISTERS[25][29] ), .ZN(n1755) );
  OAI221_X1 U1031 ( .B1(n669), .B2(n4655), .C1(n670), .C2(n4652), .A(n1763), 
        .ZN(n1760) );
  AOI22_X1 U1032 ( .A1(n4649), .A2(\REGISTERS[8][29] ), .B1(n4646), .B2(
        \REGISTERS[9][29] ), .ZN(n1763) );
  OAI221_X1 U1033 ( .B1(n619), .B2(n4703), .C1(n620), .C2(n4700), .A(n1737), 
        .ZN(n1734) );
  AOI22_X1 U1034 ( .A1(n4697), .A2(\REGISTERS[24][30] ), .B1(n4694), .B2(
        \REGISTERS[25][30] ), .ZN(n1737) );
  OAI221_X1 U1035 ( .B1(n635), .B2(n4655), .C1(n636), .C2(n4652), .A(n1745), 
        .ZN(n1742) );
  AOI22_X1 U1036 ( .A1(n4649), .A2(\REGISTERS[8][30] ), .B1(n4646), .B2(
        \REGISTERS[9][30] ), .ZN(n1745) );
  OAI221_X1 U1037 ( .B1(n558), .B2(n4703), .C1(n560), .C2(n4700), .A(n1693), 
        .ZN(n1684) );
  AOI22_X1 U1038 ( .A1(n4697), .A2(\REGISTERS[24][31] ), .B1(n4694), .B2(
        \REGISTERS[25][31] ), .ZN(n1693) );
  OAI221_X1 U1039 ( .B1(n590), .B2(n4655), .C1(n592), .C2(n4652), .A(n1717), 
        .ZN(n1708) );
  AOI22_X1 U1040 ( .A1(n4649), .A2(\REGISTERS[8][31] ), .B1(n4646), .B2(
        \REGISTERS[9][31] ), .ZN(n1717) );
  OAI221_X1 U1041 ( .B1(n4797), .B2(n1643), .C1(n4794), .C2(n1644), .A(n1645), 
        .ZN(n1634) );
  AOI22_X1 U1042 ( .A1(\REGISTERS[24][0] ), .A2(n4791), .B1(\REGISTERS[25][0] ), .B2(n4788), .ZN(n1645) );
  OAI221_X1 U1043 ( .B1(n4749), .B2(n1667), .C1(n4746), .C2(n1668), .A(n1669), 
        .ZN(n1660) );
  AOI22_X1 U1044 ( .A1(\REGISTERS[8][0] ), .A2(n4743), .B1(\REGISTERS[9][0] ), 
        .B2(n4740), .ZN(n1669) );
  OAI221_X1 U1045 ( .B1(n4797), .B2(n1605), .C1(n4794), .C2(n1606), .A(n1607), 
        .ZN(n1600) );
  AOI22_X1 U1046 ( .A1(\REGISTERS[24][1] ), .A2(n4791), .B1(\REGISTERS[25][1] ), .B2(n4788), .ZN(n1607) );
  OAI221_X1 U1047 ( .B1(n4749), .B2(n1621), .C1(n4746), .C2(n1622), .A(n1623), 
        .ZN(n1616) );
  AOI22_X1 U1048 ( .A1(\REGISTERS[8][1] ), .A2(n4743), .B1(\REGISTERS[9][1] ), 
        .B2(n4740), .ZN(n1623) );
  OAI221_X1 U1049 ( .B1(n4797), .B2(n1571), .C1(n4794), .C2(n1572), .A(n1573), 
        .ZN(n1566) );
  AOI22_X1 U1050 ( .A1(\REGISTERS[24][2] ), .A2(n4791), .B1(\REGISTERS[25][2] ), .B2(n4788), .ZN(n1573) );
  OAI221_X1 U1051 ( .B1(n4749), .B2(n1587), .C1(n4746), .C2(n1588), .A(n1589), 
        .ZN(n1582) );
  AOI22_X1 U1052 ( .A1(\REGISTERS[8][2] ), .A2(n4743), .B1(\REGISTERS[9][2] ), 
        .B2(n4740), .ZN(n1589) );
  OAI221_X1 U1053 ( .B1(n4797), .B2(n1537), .C1(n4794), .C2(n1538), .A(n1539), 
        .ZN(n1532) );
  AOI22_X1 U1054 ( .A1(\REGISTERS[24][3] ), .A2(n4791), .B1(\REGISTERS[25][3] ), .B2(n4788), .ZN(n1539) );
  OAI221_X1 U1055 ( .B1(n4749), .B2(n1553), .C1(n4746), .C2(n1554), .A(n1555), 
        .ZN(n1548) );
  AOI22_X1 U1056 ( .A1(\REGISTERS[8][3] ), .A2(n4743), .B1(\REGISTERS[9][3] ), 
        .B2(n4740), .ZN(n1555) );
  OAI221_X1 U1057 ( .B1(n4797), .B2(n1503), .C1(n4794), .C2(n1504), .A(n1505), 
        .ZN(n1498) );
  AOI22_X1 U1058 ( .A1(\REGISTERS[24][4] ), .A2(n4791), .B1(\REGISTERS[25][4] ), .B2(n4788), .ZN(n1505) );
  OAI221_X1 U1059 ( .B1(n4749), .B2(n1519), .C1(n4746), .C2(n1520), .A(n1521), 
        .ZN(n1514) );
  AOI22_X1 U1060 ( .A1(\REGISTERS[8][4] ), .A2(n4743), .B1(\REGISTERS[9][4] ), 
        .B2(n4740), .ZN(n1521) );
  OAI221_X1 U1061 ( .B1(n4797), .B2(n1469), .C1(n4794), .C2(n1470), .A(n1471), 
        .ZN(n1464) );
  AOI22_X1 U1062 ( .A1(\REGISTERS[24][5] ), .A2(n4791), .B1(\REGISTERS[25][5] ), .B2(n4788), .ZN(n1471) );
  OAI221_X1 U1063 ( .B1(n4749), .B2(n1485), .C1(n4746), .C2(n1486), .A(n1487), 
        .ZN(n1480) );
  AOI22_X1 U1064 ( .A1(\REGISTERS[8][5] ), .A2(n4743), .B1(\REGISTERS[9][5] ), 
        .B2(n4740), .ZN(n1487) );
  OAI221_X1 U1065 ( .B1(n4797), .B2(n1435), .C1(n4794), .C2(n1436), .A(n1437), 
        .ZN(n1430) );
  AOI22_X1 U1066 ( .A1(\REGISTERS[24][6] ), .A2(n4791), .B1(\REGISTERS[25][6] ), .B2(n4788), .ZN(n1437) );
  OAI221_X1 U1067 ( .B1(n4749), .B2(n1451), .C1(n4746), .C2(n1452), .A(n1453), 
        .ZN(n1446) );
  AOI22_X1 U1068 ( .A1(\REGISTERS[8][6] ), .A2(n4743), .B1(\REGISTERS[9][6] ), 
        .B2(n4740), .ZN(n1453) );
  OAI221_X1 U1069 ( .B1(n4797), .B2(n1401), .C1(n4794), .C2(n1402), .A(n1403), 
        .ZN(n1396) );
  AOI22_X1 U1070 ( .A1(\REGISTERS[24][7] ), .A2(n4791), .B1(\REGISTERS[25][7] ), .B2(n4788), .ZN(n1403) );
  OAI221_X1 U1071 ( .B1(n4749), .B2(n1417), .C1(n4746), .C2(n1418), .A(n1419), 
        .ZN(n1412) );
  AOI22_X1 U1072 ( .A1(\REGISTERS[8][7] ), .A2(n4743), .B1(\REGISTERS[9][7] ), 
        .B2(n4740), .ZN(n1419) );
  OAI221_X1 U1073 ( .B1(n4797), .B2(n1367), .C1(n4794), .C2(n1368), .A(n1369), 
        .ZN(n1362) );
  AOI22_X1 U1074 ( .A1(\REGISTERS[24][8] ), .A2(n4791), .B1(\REGISTERS[25][8] ), .B2(n4788), .ZN(n1369) );
  OAI221_X1 U1075 ( .B1(n4749), .B2(n1383), .C1(n4746), .C2(n1384), .A(n1385), 
        .ZN(n1378) );
  AOI22_X1 U1076 ( .A1(\REGISTERS[8][8] ), .A2(n4743), .B1(\REGISTERS[9][8] ), 
        .B2(n4740), .ZN(n1385) );
  OAI221_X1 U1077 ( .B1(n4797), .B2(n1333), .C1(n4794), .C2(n1334), .A(n1335), 
        .ZN(n1328) );
  AOI22_X1 U1078 ( .A1(\REGISTERS[24][9] ), .A2(n4791), .B1(\REGISTERS[25][9] ), .B2(n4788), .ZN(n1335) );
  OAI221_X1 U1079 ( .B1(n4749), .B2(n1349), .C1(n4746), .C2(n1350), .A(n1351), 
        .ZN(n1344) );
  AOI22_X1 U1080 ( .A1(\REGISTERS[8][9] ), .A2(n4743), .B1(\REGISTERS[9][9] ), 
        .B2(n4740), .ZN(n1351) );
  OAI221_X1 U1081 ( .B1(n4797), .B2(n1299), .C1(n4794), .C2(n1300), .A(n1301), 
        .ZN(n1294) );
  AOI22_X1 U1082 ( .A1(\REGISTERS[24][10] ), .A2(n4791), .B1(
        \REGISTERS[25][10] ), .B2(n4788), .ZN(n1301) );
  OAI221_X1 U1083 ( .B1(n4749), .B2(n1315), .C1(n4746), .C2(n1316), .A(n1317), 
        .ZN(n1310) );
  AOI22_X1 U1084 ( .A1(\REGISTERS[8][10] ), .A2(n4743), .B1(\REGISTERS[9][10] ), .B2(n4740), .ZN(n1317) );
  OAI221_X1 U1085 ( .B1(n4797), .B2(n1265), .C1(n4795), .C2(n1266), .A(n1267), 
        .ZN(n1260) );
  AOI22_X1 U1086 ( .A1(\REGISTERS[24][11] ), .A2(n4791), .B1(
        \REGISTERS[25][11] ), .B2(n4788), .ZN(n1267) );
  OAI221_X1 U1087 ( .B1(n4749), .B2(n1281), .C1(n4747), .C2(n1282), .A(n1283), 
        .ZN(n1276) );
  AOI22_X1 U1088 ( .A1(\REGISTERS[8][11] ), .A2(n4743), .B1(\REGISTERS[9][11] ), .B2(n4740), .ZN(n1283) );
  OAI221_X1 U1089 ( .B1(n4798), .B2(n1231), .C1(n4795), .C2(n1232), .A(n1233), 
        .ZN(n1226) );
  AOI22_X1 U1090 ( .A1(\REGISTERS[24][12] ), .A2(n4792), .B1(
        \REGISTERS[25][12] ), .B2(n4789), .ZN(n1233) );
  OAI221_X1 U1091 ( .B1(n4750), .B2(n1247), .C1(n4747), .C2(n1248), .A(n1249), 
        .ZN(n1242) );
  AOI22_X1 U1092 ( .A1(\REGISTERS[8][12] ), .A2(n4744), .B1(\REGISTERS[9][12] ), .B2(n4741), .ZN(n1249) );
  OAI221_X1 U1093 ( .B1(n4798), .B2(n1197), .C1(n4795), .C2(n1198), .A(n1199), 
        .ZN(n1192) );
  AOI22_X1 U1094 ( .A1(\REGISTERS[24][13] ), .A2(n4792), .B1(
        \REGISTERS[25][13] ), .B2(n4789), .ZN(n1199) );
  OAI221_X1 U1095 ( .B1(n4750), .B2(n1213), .C1(n4747), .C2(n1214), .A(n1215), 
        .ZN(n1208) );
  AOI22_X1 U1096 ( .A1(\REGISTERS[8][13] ), .A2(n4744), .B1(\REGISTERS[9][13] ), .B2(n4741), .ZN(n1215) );
  OAI221_X1 U1097 ( .B1(n4798), .B2(n1163), .C1(n4795), .C2(n1164), .A(n1165), 
        .ZN(n1158) );
  AOI22_X1 U1098 ( .A1(\REGISTERS[24][14] ), .A2(n4792), .B1(
        \REGISTERS[25][14] ), .B2(n4789), .ZN(n1165) );
  OAI221_X1 U1099 ( .B1(n4750), .B2(n1179), .C1(n4747), .C2(n1180), .A(n1181), 
        .ZN(n1174) );
  AOI22_X1 U1100 ( .A1(\REGISTERS[8][14] ), .A2(n4744), .B1(\REGISTERS[9][14] ), .B2(n4741), .ZN(n1181) );
  OAI221_X1 U1101 ( .B1(n4798), .B2(n1129), .C1(n4795), .C2(n1130), .A(n1131), 
        .ZN(n1124) );
  AOI22_X1 U1102 ( .A1(\REGISTERS[24][15] ), .A2(n4792), .B1(
        \REGISTERS[25][15] ), .B2(n4789), .ZN(n1131) );
  OAI221_X1 U1103 ( .B1(n4750), .B2(n1145), .C1(n4747), .C2(n1146), .A(n1147), 
        .ZN(n1140) );
  AOI22_X1 U1104 ( .A1(\REGISTERS[8][15] ), .A2(n4744), .B1(\REGISTERS[9][15] ), .B2(n4741), .ZN(n1147) );
  OAI221_X1 U1105 ( .B1(n4798), .B2(n1095), .C1(n4795), .C2(n1096), .A(n1097), 
        .ZN(n1090) );
  AOI22_X1 U1106 ( .A1(\REGISTERS[24][16] ), .A2(n4792), .B1(
        \REGISTERS[25][16] ), .B2(n4789), .ZN(n1097) );
  OAI221_X1 U1107 ( .B1(n4750), .B2(n1111), .C1(n4747), .C2(n1112), .A(n1113), 
        .ZN(n1106) );
  AOI22_X1 U1108 ( .A1(\REGISTERS[8][16] ), .A2(n4744), .B1(\REGISTERS[9][16] ), .B2(n4741), .ZN(n1113) );
  OAI221_X1 U1109 ( .B1(n4798), .B2(n1061), .C1(n4795), .C2(n1062), .A(n1063), 
        .ZN(n1056) );
  AOI22_X1 U1110 ( .A1(\REGISTERS[24][17] ), .A2(n4792), .B1(
        \REGISTERS[25][17] ), .B2(n4789), .ZN(n1063) );
  OAI221_X1 U1111 ( .B1(n4750), .B2(n1077), .C1(n4747), .C2(n1078), .A(n1079), 
        .ZN(n1072) );
  AOI22_X1 U1112 ( .A1(\REGISTERS[8][17] ), .A2(n4744), .B1(\REGISTERS[9][17] ), .B2(n4741), .ZN(n1079) );
  OAI221_X1 U1113 ( .B1(n4798), .B2(n1027), .C1(n4795), .C2(n1028), .A(n1029), 
        .ZN(n1022) );
  AOI22_X1 U1114 ( .A1(\REGISTERS[24][18] ), .A2(n4792), .B1(
        \REGISTERS[25][18] ), .B2(n4789), .ZN(n1029) );
  OAI221_X1 U1115 ( .B1(n4750), .B2(n1043), .C1(n4747), .C2(n1044), .A(n1045), 
        .ZN(n1038) );
  AOI22_X1 U1116 ( .A1(\REGISTERS[8][18] ), .A2(n4744), .B1(\REGISTERS[9][18] ), .B2(n4741), .ZN(n1045) );
  OAI221_X1 U1117 ( .B1(n4798), .B2(n993), .C1(n4795), .C2(n994), .A(n995), 
        .ZN(n988) );
  AOI22_X1 U1118 ( .A1(\REGISTERS[24][19] ), .A2(n4792), .B1(
        \REGISTERS[25][19] ), .B2(n4789), .ZN(n995) );
  OAI221_X1 U1119 ( .B1(n4750), .B2(n1009), .C1(n4747), .C2(n1010), .A(n1011), 
        .ZN(n1004) );
  AOI22_X1 U1120 ( .A1(\REGISTERS[8][19] ), .A2(n4744), .B1(\REGISTERS[9][19] ), .B2(n4741), .ZN(n1011) );
  OAI221_X1 U1121 ( .B1(n4798), .B2(n959), .C1(n4795), .C2(n960), .A(n961), 
        .ZN(n954) );
  AOI22_X1 U1122 ( .A1(\REGISTERS[24][20] ), .A2(n4792), .B1(
        \REGISTERS[25][20] ), .B2(n4789), .ZN(n961) );
  OAI221_X1 U1123 ( .B1(n4750), .B2(n975), .C1(n4747), .C2(n976), .A(n977), 
        .ZN(n970) );
  AOI22_X1 U1124 ( .A1(\REGISTERS[8][20] ), .A2(n4744), .B1(\REGISTERS[9][20] ), .B2(n4741), .ZN(n977) );
  OAI221_X1 U1125 ( .B1(n4798), .B2(n925), .C1(n4795), .C2(n926), .A(n927), 
        .ZN(n920) );
  AOI22_X1 U1126 ( .A1(\REGISTERS[24][21] ), .A2(n4792), .B1(
        \REGISTERS[25][21] ), .B2(n4789), .ZN(n927) );
  OAI221_X1 U1127 ( .B1(n4750), .B2(n941), .C1(n4747), .C2(n942), .A(n943), 
        .ZN(n936) );
  AOI22_X1 U1128 ( .A1(\REGISTERS[8][21] ), .A2(n4744), .B1(\REGISTERS[9][21] ), .B2(n4741), .ZN(n943) );
  OAI221_X1 U1129 ( .B1(n4798), .B2(n891), .C1(n4796), .C2(n892), .A(n893), 
        .ZN(n886) );
  AOI22_X1 U1130 ( .A1(\REGISTERS[24][22] ), .A2(n4792), .B1(
        \REGISTERS[25][22] ), .B2(n4789), .ZN(n893) );
  OAI221_X1 U1131 ( .B1(n4750), .B2(n907), .C1(n4748), .C2(n908), .A(n909), 
        .ZN(n902) );
  AOI22_X1 U1132 ( .A1(\REGISTERS[8][22] ), .A2(n4744), .B1(\REGISTERS[9][22] ), .B2(n4741), .ZN(n909) );
  OAI221_X1 U1133 ( .B1(n4798), .B2(n857), .C1(n4796), .C2(n858), .A(n859), 
        .ZN(n852) );
  AOI22_X1 U1134 ( .A1(\REGISTERS[24][23] ), .A2(n4792), .B1(
        \REGISTERS[25][23] ), .B2(n4789), .ZN(n859) );
  OAI221_X1 U1135 ( .B1(n4750), .B2(n873), .C1(n4748), .C2(n874), .A(n875), 
        .ZN(n868) );
  AOI22_X1 U1136 ( .A1(\REGISTERS[8][23] ), .A2(n4744), .B1(\REGISTERS[9][23] ), .B2(n4741), .ZN(n875) );
  OAI221_X1 U1137 ( .B1(n1265), .B2(n4702), .C1(n1266), .C2(n4699), .A(n2079), 
        .ZN(n2076) );
  AOI22_X1 U1138 ( .A1(n4696), .A2(\REGISTERS[24][11] ), .B1(n4693), .B2(
        \REGISTERS[25][11] ), .ZN(n2079) );
  OAI221_X1 U1139 ( .B1(n1281), .B2(n4654), .C1(n1282), .C2(n4651), .A(n2087), 
        .ZN(n2084) );
  AOI22_X1 U1140 ( .A1(n4648), .A2(\REGISTERS[8][11] ), .B1(n4645), .B2(
        \REGISTERS[9][11] ), .ZN(n2087) );
  OAI221_X1 U1141 ( .B1(n1231), .B2(n4702), .C1(n1232), .C2(n4699), .A(n2061), 
        .ZN(n2058) );
  AOI22_X1 U1142 ( .A1(n4696), .A2(\REGISTERS[24][12] ), .B1(n4693), .B2(
        \REGISTERS[25][12] ), .ZN(n2061) );
  OAI221_X1 U1143 ( .B1(n1247), .B2(n4654), .C1(n1248), .C2(n4651), .A(n2069), 
        .ZN(n2066) );
  AOI22_X1 U1144 ( .A1(n4648), .A2(\REGISTERS[8][12] ), .B1(n4645), .B2(
        \REGISTERS[9][12] ), .ZN(n2069) );
  OAI221_X1 U1145 ( .B1(n1197), .B2(n4702), .C1(n1198), .C2(n4699), .A(n2043), 
        .ZN(n2040) );
  AOI22_X1 U1146 ( .A1(n4696), .A2(\REGISTERS[24][13] ), .B1(n4693), .B2(
        \REGISTERS[25][13] ), .ZN(n2043) );
  OAI221_X1 U1147 ( .B1(n1213), .B2(n4654), .C1(n1214), .C2(n4651), .A(n2051), 
        .ZN(n2048) );
  AOI22_X1 U1148 ( .A1(n4648), .A2(\REGISTERS[8][13] ), .B1(n4645), .B2(
        \REGISTERS[9][13] ), .ZN(n2051) );
  OAI221_X1 U1149 ( .B1(n1163), .B2(n4702), .C1(n1164), .C2(n4699), .A(n2025), 
        .ZN(n2022) );
  AOI22_X1 U1150 ( .A1(n4696), .A2(\REGISTERS[24][14] ), .B1(n4693), .B2(
        \REGISTERS[25][14] ), .ZN(n2025) );
  OAI221_X1 U1151 ( .B1(n1179), .B2(n4654), .C1(n1180), .C2(n4651), .A(n2033), 
        .ZN(n2030) );
  AOI22_X1 U1152 ( .A1(n4648), .A2(\REGISTERS[8][14] ), .B1(n4645), .B2(
        \REGISTERS[9][14] ), .ZN(n2033) );
  OAI221_X1 U1153 ( .B1(n1129), .B2(n4702), .C1(n1130), .C2(n4699), .A(n2007), 
        .ZN(n2004) );
  AOI22_X1 U1154 ( .A1(n4696), .A2(\REGISTERS[24][15] ), .B1(n4693), .B2(
        \REGISTERS[25][15] ), .ZN(n2007) );
  OAI221_X1 U1155 ( .B1(n1145), .B2(n4654), .C1(n1146), .C2(n4651), .A(n2015), 
        .ZN(n2012) );
  AOI22_X1 U1156 ( .A1(n4648), .A2(\REGISTERS[8][15] ), .B1(n4645), .B2(
        \REGISTERS[9][15] ), .ZN(n2015) );
  OAI221_X1 U1157 ( .B1(n1095), .B2(n4702), .C1(n1096), .C2(n4699), .A(n1989), 
        .ZN(n1986) );
  AOI22_X1 U1158 ( .A1(n4696), .A2(\REGISTERS[24][16] ), .B1(n4693), .B2(
        \REGISTERS[25][16] ), .ZN(n1989) );
  OAI221_X1 U1159 ( .B1(n1111), .B2(n4654), .C1(n1112), .C2(n4651), .A(n1997), 
        .ZN(n1994) );
  AOI22_X1 U1160 ( .A1(n4648), .A2(\REGISTERS[8][16] ), .B1(n4645), .B2(
        \REGISTERS[9][16] ), .ZN(n1997) );
  OAI221_X1 U1161 ( .B1(n1061), .B2(n4702), .C1(n1062), .C2(n4699), .A(n1971), 
        .ZN(n1968) );
  AOI22_X1 U1162 ( .A1(n4696), .A2(\REGISTERS[24][17] ), .B1(n4693), .B2(
        \REGISTERS[25][17] ), .ZN(n1971) );
  OAI221_X1 U1163 ( .B1(n1077), .B2(n4654), .C1(n1078), .C2(n4651), .A(n1979), 
        .ZN(n1976) );
  AOI22_X1 U1164 ( .A1(n4648), .A2(\REGISTERS[8][17] ), .B1(n4645), .B2(
        \REGISTERS[9][17] ), .ZN(n1979) );
  OAI221_X1 U1165 ( .B1(n1027), .B2(n4702), .C1(n1028), .C2(n4699), .A(n1953), 
        .ZN(n1950) );
  AOI22_X1 U1166 ( .A1(n4696), .A2(\REGISTERS[24][18] ), .B1(n4693), .B2(
        \REGISTERS[25][18] ), .ZN(n1953) );
  OAI221_X1 U1167 ( .B1(n1043), .B2(n4654), .C1(n1044), .C2(n4651), .A(n1961), 
        .ZN(n1958) );
  AOI22_X1 U1168 ( .A1(n4648), .A2(\REGISTERS[8][18] ), .B1(n4645), .B2(
        \REGISTERS[9][18] ), .ZN(n1961) );
  OAI221_X1 U1169 ( .B1(n993), .B2(n4702), .C1(n994), .C2(n4699), .A(n1935), 
        .ZN(n1932) );
  AOI22_X1 U1170 ( .A1(n4696), .A2(\REGISTERS[24][19] ), .B1(n4693), .B2(
        \REGISTERS[25][19] ), .ZN(n1935) );
  OAI221_X1 U1171 ( .B1(n1009), .B2(n4654), .C1(n1010), .C2(n4651), .A(n1943), 
        .ZN(n1940) );
  AOI22_X1 U1172 ( .A1(n4648), .A2(\REGISTERS[8][19] ), .B1(n4645), .B2(
        \REGISTERS[9][19] ), .ZN(n1943) );
  OAI221_X1 U1173 ( .B1(n959), .B2(n4702), .C1(n960), .C2(n4699), .A(n1917), 
        .ZN(n1914) );
  AOI22_X1 U1174 ( .A1(n4696), .A2(\REGISTERS[24][20] ), .B1(n4693), .B2(
        \REGISTERS[25][20] ), .ZN(n1917) );
  OAI221_X1 U1175 ( .B1(n975), .B2(n4654), .C1(n976), .C2(n4651), .A(n1925), 
        .ZN(n1922) );
  AOI22_X1 U1176 ( .A1(n4648), .A2(\REGISTERS[8][20] ), .B1(n4645), .B2(
        \REGISTERS[9][20] ), .ZN(n1925) );
  OAI221_X1 U1177 ( .B1(n925), .B2(n4702), .C1(n926), .C2(n4699), .A(n1899), 
        .ZN(n1896) );
  AOI22_X1 U1178 ( .A1(n4696), .A2(\REGISTERS[24][21] ), .B1(n4693), .B2(
        \REGISTERS[25][21] ), .ZN(n1899) );
  OAI221_X1 U1179 ( .B1(n941), .B2(n4654), .C1(n942), .C2(n4651), .A(n1907), 
        .ZN(n1904) );
  AOI22_X1 U1180 ( .A1(n4648), .A2(\REGISTERS[8][21] ), .B1(n4645), .B2(
        \REGISTERS[9][21] ), .ZN(n1907) );
  OAI221_X1 U1181 ( .B1(n4787), .B2(n826), .C1(n4784), .C2(n827), .A(n828), 
        .ZN(n817) );
  AOI22_X1 U1182 ( .A1(\REGISTERS[20][24] ), .A2(n4781), .B1(
        \REGISTERS[21][24] ), .B2(n4778), .ZN(n828) );
  OAI221_X1 U1183 ( .B1(n4739), .B2(n842), .C1(n4736), .C2(n843), .A(n844), 
        .ZN(n833) );
  AOI22_X1 U1184 ( .A1(\REGISTERS[4][24] ), .A2(n4733), .B1(\REGISTERS[5][24] ), .B2(n4730), .ZN(n844) );
  OAI221_X1 U1185 ( .B1(n4787), .B2(n792), .C1(n4784), .C2(n793), .A(n794), 
        .ZN(n783) );
  AOI22_X1 U1186 ( .A1(\REGISTERS[20][25] ), .A2(n4781), .B1(
        \REGISTERS[21][25] ), .B2(n4778), .ZN(n794) );
  OAI221_X1 U1187 ( .B1(n4739), .B2(n808), .C1(n4736), .C2(n809), .A(n810), 
        .ZN(n799) );
  AOI22_X1 U1188 ( .A1(\REGISTERS[4][25] ), .A2(n4733), .B1(\REGISTERS[5][25] ), .B2(n4730), .ZN(n810) );
  OAI221_X1 U1189 ( .B1(n4787), .B2(n758), .C1(n4784), .C2(n759), .A(n760), 
        .ZN(n749) );
  AOI22_X1 U1190 ( .A1(\REGISTERS[20][26] ), .A2(n4781), .B1(
        \REGISTERS[21][26] ), .B2(n4778), .ZN(n760) );
  OAI221_X1 U1191 ( .B1(n4739), .B2(n774), .C1(n4736), .C2(n775), .A(n776), 
        .ZN(n765) );
  AOI22_X1 U1192 ( .A1(\REGISTERS[4][26] ), .A2(n4733), .B1(\REGISTERS[5][26] ), .B2(n4730), .ZN(n776) );
  OAI221_X1 U1193 ( .B1(n4787), .B2(n724), .C1(n4784), .C2(n725), .A(n726), 
        .ZN(n715) );
  AOI22_X1 U1194 ( .A1(\REGISTERS[20][27] ), .A2(n4781), .B1(
        \REGISTERS[21][27] ), .B2(n4778), .ZN(n726) );
  OAI221_X1 U1195 ( .B1(n4739), .B2(n740), .C1(n4736), .C2(n741), .A(n742), 
        .ZN(n731) );
  AOI22_X1 U1196 ( .A1(\REGISTERS[4][27] ), .A2(n4733), .B1(\REGISTERS[5][27] ), .B2(n4730), .ZN(n742) );
  OAI221_X1 U1197 ( .B1(n4787), .B2(n690), .C1(n4784), .C2(n691), .A(n692), 
        .ZN(n681) );
  AOI22_X1 U1198 ( .A1(\REGISTERS[20][28] ), .A2(n4781), .B1(
        \REGISTERS[21][28] ), .B2(n4778), .ZN(n692) );
  OAI221_X1 U1199 ( .B1(n4739), .B2(n706), .C1(n4736), .C2(n707), .A(n708), 
        .ZN(n697) );
  AOI22_X1 U1200 ( .A1(\REGISTERS[4][28] ), .A2(n4733), .B1(\REGISTERS[5][28] ), .B2(n4730), .ZN(n708) );
  OAI221_X1 U1201 ( .B1(n4787), .B2(n656), .C1(n4784), .C2(n657), .A(n658), 
        .ZN(n647) );
  AOI22_X1 U1202 ( .A1(\REGISTERS[20][29] ), .A2(n4781), .B1(
        \REGISTERS[21][29] ), .B2(n4778), .ZN(n658) );
  OAI221_X1 U1203 ( .B1(n4739), .B2(n672), .C1(n4736), .C2(n673), .A(n674), 
        .ZN(n663) );
  AOI22_X1 U1204 ( .A1(\REGISTERS[4][29] ), .A2(n4733), .B1(\REGISTERS[5][29] ), .B2(n4730), .ZN(n674) );
  OAI221_X1 U1205 ( .B1(n4787), .B2(n622), .C1(n4784), .C2(n623), .A(n624), 
        .ZN(n613) );
  AOI22_X1 U1206 ( .A1(\REGISTERS[20][30] ), .A2(n4781), .B1(
        \REGISTERS[21][30] ), .B2(n4778), .ZN(n624) );
  OAI221_X1 U1207 ( .B1(n4739), .B2(n638), .C1(n4736), .C2(n639), .A(n640), 
        .ZN(n629) );
  AOI22_X1 U1208 ( .A1(\REGISTERS[4][30] ), .A2(n4733), .B1(\REGISTERS[5][30] ), .B2(n4730), .ZN(n640) );
  OAI221_X1 U1209 ( .B1(n4787), .B2(n565), .C1(n4784), .C2(n567), .A(n568), 
        .ZN(n547) );
  AOI22_X1 U1210 ( .A1(\REGISTERS[20][31] ), .A2(n4781), .B1(
        \REGISTERS[21][31] ), .B2(n4778), .ZN(n568) );
  OAI221_X1 U1211 ( .B1(n4739), .B2(n597), .C1(n4736), .C2(n599), .A(n600), 
        .ZN(n579) );
  AOI22_X1 U1212 ( .A1(\REGISTERS[4][31] ), .A2(n4733), .B1(\REGISTERS[5][31] ), .B2(n4730), .ZN(n600) );
  OAI221_X1 U1213 ( .B1(n4775), .B2(n829), .C1(n4772), .C2(n830), .A(n831), 
        .ZN(n816) );
  AOI22_X1 U1214 ( .A1(\REGISTERS[16][24] ), .A2(n4769), .B1(
        \REGISTERS[17][24] ), .B2(n4766), .ZN(n831) );
  OAI221_X1 U1215 ( .B1(n4775), .B2(n795), .C1(n4772), .C2(n796), .A(n797), 
        .ZN(n782) );
  AOI22_X1 U1216 ( .A1(\REGISTERS[16][25] ), .A2(n4769), .B1(
        \REGISTERS[17][25] ), .B2(n4766), .ZN(n797) );
  OAI221_X1 U1217 ( .B1(n4775), .B2(n761), .C1(n4772), .C2(n762), .A(n763), 
        .ZN(n748) );
  AOI22_X1 U1218 ( .A1(\REGISTERS[16][26] ), .A2(n4769), .B1(
        \REGISTERS[17][26] ), .B2(n4766), .ZN(n763) );
  OAI221_X1 U1219 ( .B1(n4775), .B2(n727), .C1(n4772), .C2(n728), .A(n729), 
        .ZN(n714) );
  AOI22_X1 U1220 ( .A1(\REGISTERS[16][27] ), .A2(n4769), .B1(
        \REGISTERS[17][27] ), .B2(n4766), .ZN(n729) );
  OAI221_X1 U1221 ( .B1(n4775), .B2(n693), .C1(n4772), .C2(n694), .A(n695), 
        .ZN(n680) );
  AOI22_X1 U1222 ( .A1(\REGISTERS[16][28] ), .A2(n4769), .B1(
        \REGISTERS[17][28] ), .B2(n4766), .ZN(n695) );
  OAI221_X1 U1223 ( .B1(n4775), .B2(n659), .C1(n4772), .C2(n660), .A(n661), 
        .ZN(n646) );
  AOI22_X1 U1224 ( .A1(\REGISTERS[16][29] ), .A2(n4769), .B1(
        \REGISTERS[17][29] ), .B2(n4766), .ZN(n661) );
  OAI221_X1 U1225 ( .B1(n4775), .B2(n625), .C1(n4772), .C2(n626), .A(n627), 
        .ZN(n612) );
  AOI22_X1 U1226 ( .A1(\REGISTERS[16][30] ), .A2(n4769), .B1(
        \REGISTERS[17][30] ), .B2(n4766), .ZN(n627) );
  OAI221_X1 U1227 ( .B1(n4775), .B2(n572), .C1(n4772), .C2(n574), .A(n575), 
        .ZN(n546) );
  AOI22_X1 U1228 ( .A1(\REGISTERS[16][31] ), .A2(n4769), .B1(
        \REGISTERS[17][31] ), .B2(n4766), .ZN(n575) );
  OAI221_X1 U1229 ( .B1(n1649), .B2(n4689), .C1(n1650), .C2(n4686), .A(n2285), 
        .ZN(n2273) );
  AOI22_X1 U1230 ( .A1(n4683), .A2(\REGISTERS[20][0] ), .B1(n4680), .B2(
        \REGISTERS[21][0] ), .ZN(n2285) );
  OAI221_X1 U1231 ( .B1(n1670), .B2(n4641), .C1(n1671), .C2(n4638), .A(n2298), 
        .ZN(n2291) );
  AOI22_X1 U1232 ( .A1(n4635), .A2(\REGISTERS[4][0] ), .B1(n4632), .B2(
        \REGISTERS[5][0] ), .ZN(n2298) );
  OAI221_X1 U1233 ( .B1(n1608), .B2(n4689), .C1(n1609), .C2(n4686), .A(n2260), 
        .ZN(n2255) );
  AOI22_X1 U1234 ( .A1(n4683), .A2(\REGISTERS[20][1] ), .B1(n4680), .B2(
        \REGISTERS[21][1] ), .ZN(n2260) );
  OAI221_X1 U1235 ( .B1(n1624), .B2(n4641), .C1(n1625), .C2(n4638), .A(n2268), 
        .ZN(n2263) );
  AOI22_X1 U1236 ( .A1(n4635), .A2(\REGISTERS[4][1] ), .B1(n4632), .B2(
        \REGISTERS[5][1] ), .ZN(n2268) );
  OAI221_X1 U1237 ( .B1(n1574), .B2(n4689), .C1(n1575), .C2(n4686), .A(n2242), 
        .ZN(n2237) );
  AOI22_X1 U1238 ( .A1(n4683), .A2(\REGISTERS[20][2] ), .B1(n4680), .B2(
        \REGISTERS[21][2] ), .ZN(n2242) );
  OAI221_X1 U1239 ( .B1(n1590), .B2(n4641), .C1(n1591), .C2(n4638), .A(n2250), 
        .ZN(n2245) );
  AOI22_X1 U1240 ( .A1(n4635), .A2(\REGISTERS[4][2] ), .B1(n4632), .B2(
        \REGISTERS[5][2] ), .ZN(n2250) );
  OAI221_X1 U1241 ( .B1(n1540), .B2(n4689), .C1(n1541), .C2(n4686), .A(n2224), 
        .ZN(n2219) );
  AOI22_X1 U1242 ( .A1(n4683), .A2(\REGISTERS[20][3] ), .B1(n4680), .B2(
        \REGISTERS[21][3] ), .ZN(n2224) );
  OAI221_X1 U1243 ( .B1(n1556), .B2(n4641), .C1(n1557), .C2(n4638), .A(n2232), 
        .ZN(n2227) );
  AOI22_X1 U1244 ( .A1(n4635), .A2(\REGISTERS[4][3] ), .B1(n4632), .B2(
        \REGISTERS[5][3] ), .ZN(n2232) );
  OAI221_X1 U1245 ( .B1(n1506), .B2(n4689), .C1(n1507), .C2(n4686), .A(n2206), 
        .ZN(n2201) );
  AOI22_X1 U1246 ( .A1(n4683), .A2(\REGISTERS[20][4] ), .B1(n4680), .B2(
        \REGISTERS[21][4] ), .ZN(n2206) );
  OAI221_X1 U1247 ( .B1(n1522), .B2(n4641), .C1(n1523), .C2(n4638), .A(n2214), 
        .ZN(n2209) );
  AOI22_X1 U1248 ( .A1(n4635), .A2(\REGISTERS[4][4] ), .B1(n4632), .B2(
        \REGISTERS[5][4] ), .ZN(n2214) );
  OAI221_X1 U1249 ( .B1(n1472), .B2(n4689), .C1(n1473), .C2(n4686), .A(n2188), 
        .ZN(n2183) );
  AOI22_X1 U1250 ( .A1(n4683), .A2(\REGISTERS[20][5] ), .B1(n4680), .B2(
        \REGISTERS[21][5] ), .ZN(n2188) );
  OAI221_X1 U1251 ( .B1(n1488), .B2(n4641), .C1(n1489), .C2(n4638), .A(n2196), 
        .ZN(n2191) );
  AOI22_X1 U1252 ( .A1(n4635), .A2(\REGISTERS[4][5] ), .B1(n4632), .B2(
        \REGISTERS[5][5] ), .ZN(n2196) );
  OAI221_X1 U1253 ( .B1(n1438), .B2(n4689), .C1(n1439), .C2(n4686), .A(n2170), 
        .ZN(n2165) );
  AOI22_X1 U1254 ( .A1(n4683), .A2(\REGISTERS[20][6] ), .B1(n4680), .B2(
        \REGISTERS[21][6] ), .ZN(n2170) );
  OAI221_X1 U1255 ( .B1(n1454), .B2(n4641), .C1(n1455), .C2(n4638), .A(n2178), 
        .ZN(n2173) );
  AOI22_X1 U1256 ( .A1(n4635), .A2(\REGISTERS[4][6] ), .B1(n4632), .B2(
        \REGISTERS[5][6] ), .ZN(n2178) );
  OAI221_X1 U1257 ( .B1(n1404), .B2(n4689), .C1(n1405), .C2(n4686), .A(n2152), 
        .ZN(n2147) );
  AOI22_X1 U1258 ( .A1(n4683), .A2(\REGISTERS[20][7] ), .B1(n4680), .B2(
        \REGISTERS[21][7] ), .ZN(n2152) );
  OAI221_X1 U1259 ( .B1(n1420), .B2(n4641), .C1(n1421), .C2(n4638), .A(n2160), 
        .ZN(n2155) );
  AOI22_X1 U1260 ( .A1(n4635), .A2(\REGISTERS[4][7] ), .B1(n4632), .B2(
        \REGISTERS[5][7] ), .ZN(n2160) );
  OAI221_X1 U1261 ( .B1(n1370), .B2(n4689), .C1(n1371), .C2(n4686), .A(n2134), 
        .ZN(n2129) );
  AOI22_X1 U1262 ( .A1(n4683), .A2(\REGISTERS[20][8] ), .B1(n4680), .B2(
        \REGISTERS[21][8] ), .ZN(n2134) );
  OAI221_X1 U1263 ( .B1(n1386), .B2(n4641), .C1(n1387), .C2(n4638), .A(n2142), 
        .ZN(n2137) );
  AOI22_X1 U1264 ( .A1(n4635), .A2(\REGISTERS[4][8] ), .B1(n4632), .B2(
        \REGISTERS[5][8] ), .ZN(n2142) );
  OAI221_X1 U1265 ( .B1(n1336), .B2(n4689), .C1(n1337), .C2(n4686), .A(n2116), 
        .ZN(n2111) );
  AOI22_X1 U1266 ( .A1(n4683), .A2(\REGISTERS[20][9] ), .B1(n4680), .B2(
        \REGISTERS[21][9] ), .ZN(n2116) );
  OAI221_X1 U1267 ( .B1(n1352), .B2(n4641), .C1(n1353), .C2(n4638), .A(n2124), 
        .ZN(n2119) );
  AOI22_X1 U1268 ( .A1(n4635), .A2(\REGISTERS[4][9] ), .B1(n4632), .B2(
        \REGISTERS[5][9] ), .ZN(n2124) );
  OAI221_X1 U1269 ( .B1(n1302), .B2(n4689), .C1(n1303), .C2(n4686), .A(n2098), 
        .ZN(n2093) );
  AOI22_X1 U1270 ( .A1(n4683), .A2(\REGISTERS[20][10] ), .B1(n4680), .B2(
        \REGISTERS[21][10] ), .ZN(n2098) );
  OAI221_X1 U1271 ( .B1(n1318), .B2(n4641), .C1(n1319), .C2(n4638), .A(n2106), 
        .ZN(n2101) );
  AOI22_X1 U1272 ( .A1(n4635), .A2(\REGISTERS[4][10] ), .B1(n4632), .B2(
        \REGISTERS[5][10] ), .ZN(n2106) );
  OAI221_X1 U1273 ( .B1(n894), .B2(n4691), .C1(n895), .C2(n4688), .A(n1882), 
        .ZN(n1877) );
  AOI22_X1 U1274 ( .A1(n4685), .A2(\REGISTERS[20][22] ), .B1(n4682), .B2(
        \REGISTERS[21][22] ), .ZN(n1882) );
  OAI221_X1 U1275 ( .B1(n910), .B2(n4643), .C1(n911), .C2(n4640), .A(n1890), 
        .ZN(n1885) );
  AOI22_X1 U1276 ( .A1(n4637), .A2(\REGISTERS[4][22] ), .B1(n4634), .B2(
        \REGISTERS[5][22] ), .ZN(n1890) );
  OAI221_X1 U1277 ( .B1(n860), .B2(n4691), .C1(n861), .C2(n4688), .A(n1864), 
        .ZN(n1859) );
  AOI22_X1 U1278 ( .A1(n4685), .A2(\REGISTERS[20][23] ), .B1(n4682), .B2(
        \REGISTERS[21][23] ), .ZN(n1864) );
  OAI221_X1 U1279 ( .B1(n876), .B2(n4643), .C1(n877), .C2(n4640), .A(n1872), 
        .ZN(n1867) );
  AOI22_X1 U1280 ( .A1(n4637), .A2(\REGISTERS[4][23] ), .B1(n4634), .B2(
        \REGISTERS[5][23] ), .ZN(n1872) );
  OAI221_X1 U1281 ( .B1(n826), .B2(n4691), .C1(n827), .C2(n4688), .A(n1846), 
        .ZN(n1841) );
  AOI22_X1 U1282 ( .A1(n4685), .A2(\REGISTERS[20][24] ), .B1(n4682), .B2(
        \REGISTERS[21][24] ), .ZN(n1846) );
  OAI221_X1 U1283 ( .B1(n842), .B2(n4643), .C1(n843), .C2(n4640), .A(n1854), 
        .ZN(n1849) );
  AOI22_X1 U1284 ( .A1(n4637), .A2(\REGISTERS[4][24] ), .B1(n4634), .B2(
        \REGISTERS[5][24] ), .ZN(n1854) );
  OAI221_X1 U1285 ( .B1(n792), .B2(n4691), .C1(n793), .C2(n4688), .A(n1828), 
        .ZN(n1823) );
  AOI22_X1 U1286 ( .A1(n4685), .A2(\REGISTERS[20][25] ), .B1(n4682), .B2(
        \REGISTERS[21][25] ), .ZN(n1828) );
  OAI221_X1 U1287 ( .B1(n808), .B2(n4643), .C1(n809), .C2(n4640), .A(n1836), 
        .ZN(n1831) );
  AOI22_X1 U1288 ( .A1(n4637), .A2(\REGISTERS[4][25] ), .B1(n4634), .B2(
        \REGISTERS[5][25] ), .ZN(n1836) );
  OAI221_X1 U1289 ( .B1(n758), .B2(n4691), .C1(n759), .C2(n4688), .A(n1810), 
        .ZN(n1805) );
  AOI22_X1 U1290 ( .A1(n4685), .A2(\REGISTERS[20][26] ), .B1(n4682), .B2(
        \REGISTERS[21][26] ), .ZN(n1810) );
  OAI221_X1 U1291 ( .B1(n774), .B2(n4643), .C1(n775), .C2(n4640), .A(n1818), 
        .ZN(n1813) );
  AOI22_X1 U1292 ( .A1(n4637), .A2(\REGISTERS[4][26] ), .B1(n4634), .B2(
        \REGISTERS[5][26] ), .ZN(n1818) );
  OAI221_X1 U1293 ( .B1(n724), .B2(n4691), .C1(n725), .C2(n4688), .A(n1792), 
        .ZN(n1787) );
  AOI22_X1 U1294 ( .A1(n4685), .A2(\REGISTERS[20][27] ), .B1(n4682), .B2(
        \REGISTERS[21][27] ), .ZN(n1792) );
  OAI221_X1 U1295 ( .B1(n740), .B2(n4643), .C1(n741), .C2(n4640), .A(n1800), 
        .ZN(n1795) );
  AOI22_X1 U1296 ( .A1(n4637), .A2(\REGISTERS[4][27] ), .B1(n4634), .B2(
        \REGISTERS[5][27] ), .ZN(n1800) );
  OAI221_X1 U1297 ( .B1(n690), .B2(n4691), .C1(n691), .C2(n4688), .A(n1774), 
        .ZN(n1769) );
  AOI22_X1 U1298 ( .A1(n4685), .A2(\REGISTERS[20][28] ), .B1(n4682), .B2(
        \REGISTERS[21][28] ), .ZN(n1774) );
  OAI221_X1 U1299 ( .B1(n706), .B2(n4643), .C1(n707), .C2(n4640), .A(n1782), 
        .ZN(n1777) );
  AOI22_X1 U1300 ( .A1(n4637), .A2(\REGISTERS[4][28] ), .B1(n4634), .B2(
        \REGISTERS[5][28] ), .ZN(n1782) );
  OAI221_X1 U1301 ( .B1(n656), .B2(n4691), .C1(n657), .C2(n4688), .A(n1756), 
        .ZN(n1751) );
  AOI22_X1 U1302 ( .A1(n4685), .A2(\REGISTERS[20][29] ), .B1(n4682), .B2(
        \REGISTERS[21][29] ), .ZN(n1756) );
  OAI221_X1 U1303 ( .B1(n672), .B2(n4643), .C1(n673), .C2(n4640), .A(n1764), 
        .ZN(n1759) );
  AOI22_X1 U1304 ( .A1(n4637), .A2(\REGISTERS[4][29] ), .B1(n4634), .B2(
        \REGISTERS[5][29] ), .ZN(n1764) );
  OAI221_X1 U1305 ( .B1(n622), .B2(n4691), .C1(n623), .C2(n4688), .A(n1738), 
        .ZN(n1733) );
  AOI22_X1 U1306 ( .A1(n4685), .A2(\REGISTERS[20][30] ), .B1(n4682), .B2(
        \REGISTERS[21][30] ), .ZN(n1738) );
  OAI221_X1 U1307 ( .B1(n638), .B2(n4643), .C1(n639), .C2(n4640), .A(n1746), 
        .ZN(n1741) );
  AOI22_X1 U1308 ( .A1(n4637), .A2(\REGISTERS[4][30] ), .B1(n4634), .B2(
        \REGISTERS[5][30] ), .ZN(n1746) );
  OAI221_X1 U1309 ( .B1(n565), .B2(n4691), .C1(n567), .C2(n4688), .A(n1698), 
        .ZN(n1683) );
  AOI22_X1 U1310 ( .A1(n4685), .A2(\REGISTERS[20][31] ), .B1(n4682), .B2(
        \REGISTERS[21][31] ), .ZN(n1698) );
  OAI221_X1 U1311 ( .B1(n597), .B2(n4643), .C1(n599), .C2(n4640), .A(n1722), 
        .ZN(n1707) );
  AOI22_X1 U1312 ( .A1(n4637), .A2(\REGISTERS[4][31] ), .B1(n4634), .B2(
        \REGISTERS[5][31] ), .ZN(n1722) );
  OAI221_X1 U1313 ( .B1(n1654), .B2(n4677), .C1(n1655), .C2(n4674), .A(n2288), 
        .ZN(n2272) );
  AOI22_X1 U1314 ( .A1(n4671), .A2(\REGISTERS[16][0] ), .B1(n4668), .B2(
        \REGISTERS[17][0] ), .ZN(n2288) );
  OAI221_X1 U1315 ( .B1(n1611), .B2(n4677), .C1(n1612), .C2(n4674), .A(n2261), 
        .ZN(n2254) );
  AOI22_X1 U1316 ( .A1(n4671), .A2(\REGISTERS[16][1] ), .B1(n4668), .B2(
        \REGISTERS[17][1] ), .ZN(n2261) );
  OAI221_X1 U1317 ( .B1(n1577), .B2(n4677), .C1(n1578), .C2(n4674), .A(n2243), 
        .ZN(n2236) );
  AOI22_X1 U1318 ( .A1(n4671), .A2(\REGISTERS[16][2] ), .B1(n4668), .B2(
        \REGISTERS[17][2] ), .ZN(n2243) );
  OAI221_X1 U1319 ( .B1(n1543), .B2(n4677), .C1(n1544), .C2(n4674), .A(n2225), 
        .ZN(n2218) );
  AOI22_X1 U1320 ( .A1(n4671), .A2(\REGISTERS[16][3] ), .B1(n4668), .B2(
        \REGISTERS[17][3] ), .ZN(n2225) );
  OAI221_X1 U1321 ( .B1(n1509), .B2(n4677), .C1(n1510), .C2(n4674), .A(n2207), 
        .ZN(n2200) );
  AOI22_X1 U1322 ( .A1(n4671), .A2(\REGISTERS[16][4] ), .B1(n4668), .B2(
        \REGISTERS[17][4] ), .ZN(n2207) );
  OAI221_X1 U1323 ( .B1(n1475), .B2(n4677), .C1(n1476), .C2(n4674), .A(n2189), 
        .ZN(n2182) );
  AOI22_X1 U1324 ( .A1(n4671), .A2(\REGISTERS[16][5] ), .B1(n4668), .B2(
        \REGISTERS[17][5] ), .ZN(n2189) );
  OAI221_X1 U1325 ( .B1(n1441), .B2(n4677), .C1(n1442), .C2(n4674), .A(n2171), 
        .ZN(n2164) );
  AOI22_X1 U1326 ( .A1(n4671), .A2(\REGISTERS[16][6] ), .B1(n4668), .B2(
        \REGISTERS[17][6] ), .ZN(n2171) );
  OAI221_X1 U1327 ( .B1(n1407), .B2(n4677), .C1(n1408), .C2(n4674), .A(n2153), 
        .ZN(n2146) );
  AOI22_X1 U1328 ( .A1(n4671), .A2(\REGISTERS[16][7] ), .B1(n4668), .B2(
        \REGISTERS[17][7] ), .ZN(n2153) );
  OAI221_X1 U1329 ( .B1(n1373), .B2(n4677), .C1(n1374), .C2(n4674), .A(n2135), 
        .ZN(n2128) );
  AOI22_X1 U1330 ( .A1(n4671), .A2(\REGISTERS[16][8] ), .B1(n4668), .B2(
        \REGISTERS[17][8] ), .ZN(n2135) );
  OAI221_X1 U1331 ( .B1(n1339), .B2(n4677), .C1(n1340), .C2(n4674), .A(n2117), 
        .ZN(n2110) );
  AOI22_X1 U1332 ( .A1(n4671), .A2(\REGISTERS[16][9] ), .B1(n4668), .B2(
        \REGISTERS[17][9] ), .ZN(n2117) );
  OAI221_X1 U1333 ( .B1(n1305), .B2(n4677), .C1(n1306), .C2(n4674), .A(n2099), 
        .ZN(n2092) );
  AOI22_X1 U1334 ( .A1(n4671), .A2(\REGISTERS[16][10] ), .B1(n4668), .B2(
        \REGISTERS[17][10] ), .ZN(n2099) );
  OAI221_X1 U1335 ( .B1(n897), .B2(n4679), .C1(n898), .C2(n4676), .A(n1883), 
        .ZN(n1876) );
  AOI22_X1 U1336 ( .A1(n4673), .A2(\REGISTERS[16][22] ), .B1(n4670), .B2(
        \REGISTERS[17][22] ), .ZN(n1883) );
  OAI221_X1 U1337 ( .B1(n863), .B2(n4679), .C1(n864), .C2(n4676), .A(n1865), 
        .ZN(n1858) );
  AOI22_X1 U1338 ( .A1(n4673), .A2(\REGISTERS[16][23] ), .B1(n4670), .B2(
        \REGISTERS[17][23] ), .ZN(n1865) );
  OAI221_X1 U1339 ( .B1(n829), .B2(n4679), .C1(n830), .C2(n4676), .A(n1847), 
        .ZN(n1840) );
  AOI22_X1 U1340 ( .A1(n4673), .A2(\REGISTERS[16][24] ), .B1(n4670), .B2(
        \REGISTERS[17][24] ), .ZN(n1847) );
  OAI221_X1 U1341 ( .B1(n795), .B2(n4679), .C1(n796), .C2(n4676), .A(n1829), 
        .ZN(n1822) );
  AOI22_X1 U1342 ( .A1(n4673), .A2(\REGISTERS[16][25] ), .B1(n4670), .B2(
        \REGISTERS[17][25] ), .ZN(n1829) );
  OAI221_X1 U1343 ( .B1(n761), .B2(n4679), .C1(n762), .C2(n4676), .A(n1811), 
        .ZN(n1804) );
  AOI22_X1 U1344 ( .A1(n4673), .A2(\REGISTERS[16][26] ), .B1(n4670), .B2(
        \REGISTERS[17][26] ), .ZN(n1811) );
  OAI221_X1 U1345 ( .B1(n727), .B2(n4679), .C1(n728), .C2(n4676), .A(n1793), 
        .ZN(n1786) );
  AOI22_X1 U1346 ( .A1(n4673), .A2(\REGISTERS[16][27] ), .B1(n4670), .B2(
        \REGISTERS[17][27] ), .ZN(n1793) );
  OAI221_X1 U1347 ( .B1(n693), .B2(n4679), .C1(n694), .C2(n4676), .A(n1775), 
        .ZN(n1768) );
  AOI22_X1 U1348 ( .A1(n4673), .A2(\REGISTERS[16][28] ), .B1(n4670), .B2(
        \REGISTERS[17][28] ), .ZN(n1775) );
  OAI221_X1 U1349 ( .B1(n659), .B2(n4679), .C1(n660), .C2(n4676), .A(n1757), 
        .ZN(n1750) );
  AOI22_X1 U1350 ( .A1(n4673), .A2(\REGISTERS[16][29] ), .B1(n4670), .B2(
        \REGISTERS[17][29] ), .ZN(n1757) );
  OAI221_X1 U1351 ( .B1(n625), .B2(n4679), .C1(n626), .C2(n4676), .A(n1739), 
        .ZN(n1732) );
  AOI22_X1 U1352 ( .A1(n4673), .A2(\REGISTERS[16][30] ), .B1(n4670), .B2(
        \REGISTERS[17][30] ), .ZN(n1739) );
  OAI221_X1 U1353 ( .B1(n572), .B2(n4679), .C1(n574), .C2(n4676), .A(n1703), 
        .ZN(n1682) );
  AOI22_X1 U1354 ( .A1(n4673), .A2(\REGISTERS[16][31] ), .B1(n4670), .B2(
        \REGISTERS[17][31] ), .ZN(n1703) );
  OAI221_X1 U1355 ( .B1(n4785), .B2(n1649), .C1(n4782), .C2(n1650), .A(n1651), 
        .ZN(n1633) );
  AOI22_X1 U1356 ( .A1(\REGISTERS[20][0] ), .A2(n4779), .B1(\REGISTERS[21][0] ), .B2(n4776), .ZN(n1651) );
  OAI221_X1 U1357 ( .B1(n4737), .B2(n1670), .C1(n4734), .C2(n1671), .A(n1672), 
        .ZN(n1659) );
  AOI22_X1 U1358 ( .A1(\REGISTERS[4][0] ), .A2(n4731), .B1(\REGISTERS[5][0] ), 
        .B2(n4728), .ZN(n1672) );
  OAI221_X1 U1359 ( .B1(n4785), .B2(n1608), .C1(n4782), .C2(n1609), .A(n1610), 
        .ZN(n1599) );
  AOI22_X1 U1360 ( .A1(\REGISTERS[20][1] ), .A2(n4779), .B1(\REGISTERS[21][1] ), .B2(n4776), .ZN(n1610) );
  OAI221_X1 U1361 ( .B1(n4737), .B2(n1624), .C1(n4734), .C2(n1625), .A(n1626), 
        .ZN(n1615) );
  AOI22_X1 U1362 ( .A1(\REGISTERS[4][1] ), .A2(n4731), .B1(\REGISTERS[5][1] ), 
        .B2(n4728), .ZN(n1626) );
  OAI221_X1 U1363 ( .B1(n4785), .B2(n1574), .C1(n4782), .C2(n1575), .A(n1576), 
        .ZN(n1565) );
  AOI22_X1 U1364 ( .A1(\REGISTERS[20][2] ), .A2(n4779), .B1(\REGISTERS[21][2] ), .B2(n4776), .ZN(n1576) );
  OAI221_X1 U1365 ( .B1(n4737), .B2(n1590), .C1(n4734), .C2(n1591), .A(n1592), 
        .ZN(n1581) );
  AOI22_X1 U1366 ( .A1(\REGISTERS[4][2] ), .A2(n4731), .B1(\REGISTERS[5][2] ), 
        .B2(n4728), .ZN(n1592) );
  OAI221_X1 U1367 ( .B1(n4785), .B2(n1540), .C1(n4782), .C2(n1541), .A(n1542), 
        .ZN(n1531) );
  AOI22_X1 U1368 ( .A1(\REGISTERS[20][3] ), .A2(n4779), .B1(\REGISTERS[21][3] ), .B2(n4776), .ZN(n1542) );
  OAI221_X1 U1369 ( .B1(n4737), .B2(n1556), .C1(n4734), .C2(n1557), .A(n1558), 
        .ZN(n1547) );
  AOI22_X1 U1370 ( .A1(\REGISTERS[4][3] ), .A2(n4731), .B1(\REGISTERS[5][3] ), 
        .B2(n4728), .ZN(n1558) );
  OAI221_X1 U1371 ( .B1(n4785), .B2(n1506), .C1(n4782), .C2(n1507), .A(n1508), 
        .ZN(n1497) );
  AOI22_X1 U1372 ( .A1(\REGISTERS[20][4] ), .A2(n4779), .B1(\REGISTERS[21][4] ), .B2(n4776), .ZN(n1508) );
  OAI221_X1 U1373 ( .B1(n4737), .B2(n1522), .C1(n4734), .C2(n1523), .A(n1524), 
        .ZN(n1513) );
  AOI22_X1 U1374 ( .A1(\REGISTERS[4][4] ), .A2(n4731), .B1(\REGISTERS[5][4] ), 
        .B2(n4728), .ZN(n1524) );
  OAI221_X1 U1375 ( .B1(n4785), .B2(n1472), .C1(n4782), .C2(n1473), .A(n1474), 
        .ZN(n1463) );
  AOI22_X1 U1376 ( .A1(\REGISTERS[20][5] ), .A2(n4779), .B1(\REGISTERS[21][5] ), .B2(n4776), .ZN(n1474) );
  OAI221_X1 U1377 ( .B1(n4737), .B2(n1488), .C1(n4734), .C2(n1489), .A(n1490), 
        .ZN(n1479) );
  AOI22_X1 U1378 ( .A1(\REGISTERS[4][5] ), .A2(n4731), .B1(\REGISTERS[5][5] ), 
        .B2(n4728), .ZN(n1490) );
  OAI221_X1 U1379 ( .B1(n4785), .B2(n1438), .C1(n4782), .C2(n1439), .A(n1440), 
        .ZN(n1429) );
  AOI22_X1 U1380 ( .A1(\REGISTERS[20][6] ), .A2(n4779), .B1(\REGISTERS[21][6] ), .B2(n4776), .ZN(n1440) );
  OAI221_X1 U1381 ( .B1(n4737), .B2(n1454), .C1(n4734), .C2(n1455), .A(n1456), 
        .ZN(n1445) );
  AOI22_X1 U1382 ( .A1(\REGISTERS[4][6] ), .A2(n4731), .B1(\REGISTERS[5][6] ), 
        .B2(n4728), .ZN(n1456) );
  OAI221_X1 U1383 ( .B1(n4785), .B2(n1404), .C1(n4782), .C2(n1405), .A(n1406), 
        .ZN(n1395) );
  AOI22_X1 U1384 ( .A1(\REGISTERS[20][7] ), .A2(n4779), .B1(\REGISTERS[21][7] ), .B2(n4776), .ZN(n1406) );
  OAI221_X1 U1385 ( .B1(n4737), .B2(n1420), .C1(n4734), .C2(n1421), .A(n1422), 
        .ZN(n1411) );
  AOI22_X1 U1386 ( .A1(\REGISTERS[4][7] ), .A2(n4731), .B1(\REGISTERS[5][7] ), 
        .B2(n4728), .ZN(n1422) );
  OAI221_X1 U1387 ( .B1(n4785), .B2(n1370), .C1(n4782), .C2(n1371), .A(n1372), 
        .ZN(n1361) );
  AOI22_X1 U1388 ( .A1(\REGISTERS[20][8] ), .A2(n4779), .B1(\REGISTERS[21][8] ), .B2(n4776), .ZN(n1372) );
  OAI221_X1 U1389 ( .B1(n4737), .B2(n1386), .C1(n4734), .C2(n1387), .A(n1388), 
        .ZN(n1377) );
  AOI22_X1 U1390 ( .A1(\REGISTERS[4][8] ), .A2(n4731), .B1(\REGISTERS[5][8] ), 
        .B2(n4728), .ZN(n1388) );
  OAI221_X1 U1391 ( .B1(n4785), .B2(n1336), .C1(n4782), .C2(n1337), .A(n1338), 
        .ZN(n1327) );
  AOI22_X1 U1392 ( .A1(\REGISTERS[20][9] ), .A2(n4779), .B1(\REGISTERS[21][9] ), .B2(n4776), .ZN(n1338) );
  OAI221_X1 U1393 ( .B1(n4737), .B2(n1352), .C1(n4734), .C2(n1353), .A(n1354), 
        .ZN(n1343) );
  AOI22_X1 U1394 ( .A1(\REGISTERS[4][9] ), .A2(n4731), .B1(\REGISTERS[5][9] ), 
        .B2(n4728), .ZN(n1354) );
  OAI221_X1 U1395 ( .B1(n4785), .B2(n1302), .C1(n4782), .C2(n1303), .A(n1304), 
        .ZN(n1293) );
  AOI22_X1 U1396 ( .A1(\REGISTERS[20][10] ), .A2(n4779), .B1(
        \REGISTERS[21][10] ), .B2(n4776), .ZN(n1304) );
  OAI221_X1 U1397 ( .B1(n4737), .B2(n1318), .C1(n4734), .C2(n1319), .A(n1320), 
        .ZN(n1309) );
  AOI22_X1 U1398 ( .A1(\REGISTERS[4][10] ), .A2(n4731), .B1(\REGISTERS[5][10] ), .B2(n4728), .ZN(n1320) );
  OAI221_X1 U1399 ( .B1(n4785), .B2(n1268), .C1(n4783), .C2(n1269), .A(n1270), 
        .ZN(n1259) );
  AOI22_X1 U1400 ( .A1(\REGISTERS[20][11] ), .A2(n4779), .B1(
        \REGISTERS[21][11] ), .B2(n4776), .ZN(n1270) );
  OAI221_X1 U1401 ( .B1(n4737), .B2(n1284), .C1(n4735), .C2(n1285), .A(n1286), 
        .ZN(n1275) );
  AOI22_X1 U1402 ( .A1(\REGISTERS[4][11] ), .A2(n4731), .B1(\REGISTERS[5][11] ), .B2(n4728), .ZN(n1286) );
  OAI221_X1 U1403 ( .B1(n4786), .B2(n1234), .C1(n4783), .C2(n1235), .A(n1236), 
        .ZN(n1225) );
  AOI22_X1 U1404 ( .A1(\REGISTERS[20][12] ), .A2(n4780), .B1(
        \REGISTERS[21][12] ), .B2(n4777), .ZN(n1236) );
  OAI221_X1 U1405 ( .B1(n4738), .B2(n1250), .C1(n4735), .C2(n1251), .A(n1252), 
        .ZN(n1241) );
  AOI22_X1 U1406 ( .A1(\REGISTERS[4][12] ), .A2(n4732), .B1(\REGISTERS[5][12] ), .B2(n4729), .ZN(n1252) );
  OAI221_X1 U1407 ( .B1(n4786), .B2(n1200), .C1(n4783), .C2(n1201), .A(n1202), 
        .ZN(n1191) );
  AOI22_X1 U1408 ( .A1(\REGISTERS[20][13] ), .A2(n4780), .B1(
        \REGISTERS[21][13] ), .B2(n4777), .ZN(n1202) );
  OAI221_X1 U1409 ( .B1(n4738), .B2(n1216), .C1(n4735), .C2(n1217), .A(n1218), 
        .ZN(n1207) );
  AOI22_X1 U1410 ( .A1(\REGISTERS[4][13] ), .A2(n4732), .B1(\REGISTERS[5][13] ), .B2(n4729), .ZN(n1218) );
  OAI221_X1 U1411 ( .B1(n4786), .B2(n1166), .C1(n4783), .C2(n1167), .A(n1168), 
        .ZN(n1157) );
  AOI22_X1 U1412 ( .A1(\REGISTERS[20][14] ), .A2(n4780), .B1(
        \REGISTERS[21][14] ), .B2(n4777), .ZN(n1168) );
  OAI221_X1 U1413 ( .B1(n4738), .B2(n1182), .C1(n4735), .C2(n1183), .A(n1184), 
        .ZN(n1173) );
  AOI22_X1 U1414 ( .A1(\REGISTERS[4][14] ), .A2(n4732), .B1(\REGISTERS[5][14] ), .B2(n4729), .ZN(n1184) );
  OAI221_X1 U1415 ( .B1(n4786), .B2(n1132), .C1(n4783), .C2(n1133), .A(n1134), 
        .ZN(n1123) );
  AOI22_X1 U1416 ( .A1(\REGISTERS[20][15] ), .A2(n4780), .B1(
        \REGISTERS[21][15] ), .B2(n4777), .ZN(n1134) );
  OAI221_X1 U1417 ( .B1(n4738), .B2(n1148), .C1(n4735), .C2(n1149), .A(n1150), 
        .ZN(n1139) );
  AOI22_X1 U1418 ( .A1(\REGISTERS[4][15] ), .A2(n4732), .B1(\REGISTERS[5][15] ), .B2(n4729), .ZN(n1150) );
  OAI221_X1 U1419 ( .B1(n4786), .B2(n1098), .C1(n4783), .C2(n1099), .A(n1100), 
        .ZN(n1089) );
  AOI22_X1 U1420 ( .A1(\REGISTERS[20][16] ), .A2(n4780), .B1(
        \REGISTERS[21][16] ), .B2(n4777), .ZN(n1100) );
  OAI221_X1 U1421 ( .B1(n4738), .B2(n1114), .C1(n4735), .C2(n1115), .A(n1116), 
        .ZN(n1105) );
  AOI22_X1 U1422 ( .A1(\REGISTERS[4][16] ), .A2(n4732), .B1(\REGISTERS[5][16] ), .B2(n4729), .ZN(n1116) );
  OAI221_X1 U1423 ( .B1(n4786), .B2(n1064), .C1(n4783), .C2(n1065), .A(n1066), 
        .ZN(n1055) );
  AOI22_X1 U1424 ( .A1(\REGISTERS[20][17] ), .A2(n4780), .B1(
        \REGISTERS[21][17] ), .B2(n4777), .ZN(n1066) );
  OAI221_X1 U1425 ( .B1(n4738), .B2(n1080), .C1(n4735), .C2(n1081), .A(n1082), 
        .ZN(n1071) );
  AOI22_X1 U1426 ( .A1(\REGISTERS[4][17] ), .A2(n4732), .B1(\REGISTERS[5][17] ), .B2(n4729), .ZN(n1082) );
  OAI221_X1 U1427 ( .B1(n4786), .B2(n1030), .C1(n4783), .C2(n1031), .A(n1032), 
        .ZN(n1021) );
  AOI22_X1 U1428 ( .A1(\REGISTERS[20][18] ), .A2(n4780), .B1(
        \REGISTERS[21][18] ), .B2(n4777), .ZN(n1032) );
  OAI221_X1 U1429 ( .B1(n4738), .B2(n1046), .C1(n4735), .C2(n1047), .A(n1048), 
        .ZN(n1037) );
  AOI22_X1 U1430 ( .A1(\REGISTERS[4][18] ), .A2(n4732), .B1(\REGISTERS[5][18] ), .B2(n4729), .ZN(n1048) );
  OAI221_X1 U1431 ( .B1(n4786), .B2(n996), .C1(n4783), .C2(n997), .A(n998), 
        .ZN(n987) );
  AOI22_X1 U1432 ( .A1(\REGISTERS[20][19] ), .A2(n4780), .B1(
        \REGISTERS[21][19] ), .B2(n4777), .ZN(n998) );
  OAI221_X1 U1433 ( .B1(n4738), .B2(n1012), .C1(n4735), .C2(n1013), .A(n1014), 
        .ZN(n1003) );
  AOI22_X1 U1434 ( .A1(\REGISTERS[4][19] ), .A2(n4732), .B1(\REGISTERS[5][19] ), .B2(n4729), .ZN(n1014) );
  OAI221_X1 U1435 ( .B1(n4786), .B2(n962), .C1(n4783), .C2(n963), .A(n964), 
        .ZN(n953) );
  AOI22_X1 U1436 ( .A1(\REGISTERS[20][20] ), .A2(n4780), .B1(
        \REGISTERS[21][20] ), .B2(n4777), .ZN(n964) );
  OAI221_X1 U1437 ( .B1(n4738), .B2(n978), .C1(n4735), .C2(n979), .A(n980), 
        .ZN(n969) );
  AOI22_X1 U1438 ( .A1(\REGISTERS[4][20] ), .A2(n4732), .B1(\REGISTERS[5][20] ), .B2(n4729), .ZN(n980) );
  OAI221_X1 U1439 ( .B1(n4786), .B2(n928), .C1(n4783), .C2(n929), .A(n930), 
        .ZN(n919) );
  AOI22_X1 U1440 ( .A1(\REGISTERS[20][21] ), .A2(n4780), .B1(
        \REGISTERS[21][21] ), .B2(n4777), .ZN(n930) );
  OAI221_X1 U1441 ( .B1(n4738), .B2(n944), .C1(n4735), .C2(n945), .A(n946), 
        .ZN(n935) );
  AOI22_X1 U1442 ( .A1(\REGISTERS[4][21] ), .A2(n4732), .B1(\REGISTERS[5][21] ), .B2(n4729), .ZN(n946) );
  OAI221_X1 U1443 ( .B1(n4786), .B2(n894), .C1(n4784), .C2(n895), .A(n896), 
        .ZN(n885) );
  AOI22_X1 U1444 ( .A1(\REGISTERS[20][22] ), .A2(n4780), .B1(
        \REGISTERS[21][22] ), .B2(n4777), .ZN(n896) );
  OAI221_X1 U1445 ( .B1(n4738), .B2(n910), .C1(n4736), .C2(n911), .A(n912), 
        .ZN(n901) );
  AOI22_X1 U1446 ( .A1(\REGISTERS[4][22] ), .A2(n4732), .B1(\REGISTERS[5][22] ), .B2(n4729), .ZN(n912) );
  OAI221_X1 U1447 ( .B1(n4786), .B2(n860), .C1(n4784), .C2(n861), .A(n862), 
        .ZN(n851) );
  AOI22_X1 U1448 ( .A1(\REGISTERS[20][23] ), .A2(n4780), .B1(
        \REGISTERS[21][23] ), .B2(n4777), .ZN(n862) );
  OAI221_X1 U1449 ( .B1(n4738), .B2(n876), .C1(n4736), .C2(n877), .A(n878), 
        .ZN(n867) );
  AOI22_X1 U1450 ( .A1(\REGISTERS[4][23] ), .A2(n4732), .B1(\REGISTERS[5][23] ), .B2(n4729), .ZN(n878) );
  OAI221_X1 U1451 ( .B1(n1268), .B2(n4690), .C1(n1269), .C2(n4687), .A(n2080), 
        .ZN(n2075) );
  AOI22_X1 U1452 ( .A1(n4684), .A2(\REGISTERS[20][11] ), .B1(n4681), .B2(
        \REGISTERS[21][11] ), .ZN(n2080) );
  OAI221_X1 U1453 ( .B1(n1284), .B2(n4642), .C1(n1285), .C2(n4639), .A(n2088), 
        .ZN(n2083) );
  AOI22_X1 U1454 ( .A1(n4636), .A2(\REGISTERS[4][11] ), .B1(n4633), .B2(
        \REGISTERS[5][11] ), .ZN(n2088) );
  OAI221_X1 U1455 ( .B1(n1234), .B2(n4690), .C1(n1235), .C2(n4687), .A(n2062), 
        .ZN(n2057) );
  AOI22_X1 U1456 ( .A1(n4684), .A2(\REGISTERS[20][12] ), .B1(n4681), .B2(
        \REGISTERS[21][12] ), .ZN(n2062) );
  OAI221_X1 U1457 ( .B1(n1250), .B2(n4642), .C1(n1251), .C2(n4639), .A(n2070), 
        .ZN(n2065) );
  AOI22_X1 U1458 ( .A1(n4636), .A2(\REGISTERS[4][12] ), .B1(n4633), .B2(
        \REGISTERS[5][12] ), .ZN(n2070) );
  OAI221_X1 U1459 ( .B1(n1200), .B2(n4690), .C1(n1201), .C2(n4687), .A(n2044), 
        .ZN(n2039) );
  AOI22_X1 U1460 ( .A1(n4684), .A2(\REGISTERS[20][13] ), .B1(n4681), .B2(
        \REGISTERS[21][13] ), .ZN(n2044) );
  OAI221_X1 U1461 ( .B1(n1216), .B2(n4642), .C1(n1217), .C2(n4639), .A(n2052), 
        .ZN(n2047) );
  AOI22_X1 U1462 ( .A1(n4636), .A2(\REGISTERS[4][13] ), .B1(n4633), .B2(
        \REGISTERS[5][13] ), .ZN(n2052) );
  OAI221_X1 U1463 ( .B1(n1166), .B2(n4690), .C1(n1167), .C2(n4687), .A(n2026), 
        .ZN(n2021) );
  AOI22_X1 U1464 ( .A1(n4684), .A2(\REGISTERS[20][14] ), .B1(n4681), .B2(
        \REGISTERS[21][14] ), .ZN(n2026) );
  OAI221_X1 U1465 ( .B1(n1182), .B2(n4642), .C1(n1183), .C2(n4639), .A(n2034), 
        .ZN(n2029) );
  AOI22_X1 U1466 ( .A1(n4636), .A2(\REGISTERS[4][14] ), .B1(n4633), .B2(
        \REGISTERS[5][14] ), .ZN(n2034) );
  OAI221_X1 U1467 ( .B1(n1132), .B2(n4690), .C1(n1133), .C2(n4687), .A(n2008), 
        .ZN(n2003) );
  AOI22_X1 U1468 ( .A1(n4684), .A2(\REGISTERS[20][15] ), .B1(n4681), .B2(
        \REGISTERS[21][15] ), .ZN(n2008) );
  OAI221_X1 U1469 ( .B1(n1148), .B2(n4642), .C1(n1149), .C2(n4639), .A(n2016), 
        .ZN(n2011) );
  AOI22_X1 U1470 ( .A1(n4636), .A2(\REGISTERS[4][15] ), .B1(n4633), .B2(
        \REGISTERS[5][15] ), .ZN(n2016) );
  OAI221_X1 U1471 ( .B1(n1098), .B2(n4690), .C1(n1099), .C2(n4687), .A(n1990), 
        .ZN(n1985) );
  AOI22_X1 U1472 ( .A1(n4684), .A2(\REGISTERS[20][16] ), .B1(n4681), .B2(
        \REGISTERS[21][16] ), .ZN(n1990) );
  OAI221_X1 U1473 ( .B1(n1114), .B2(n4642), .C1(n1115), .C2(n4639), .A(n1998), 
        .ZN(n1993) );
  AOI22_X1 U1474 ( .A1(n4636), .A2(\REGISTERS[4][16] ), .B1(n4633), .B2(
        \REGISTERS[5][16] ), .ZN(n1998) );
  OAI221_X1 U1475 ( .B1(n1064), .B2(n4690), .C1(n1065), .C2(n4687), .A(n1972), 
        .ZN(n1967) );
  AOI22_X1 U1476 ( .A1(n4684), .A2(\REGISTERS[20][17] ), .B1(n4681), .B2(
        \REGISTERS[21][17] ), .ZN(n1972) );
  OAI221_X1 U1477 ( .B1(n1080), .B2(n4642), .C1(n1081), .C2(n4639), .A(n1980), 
        .ZN(n1975) );
  AOI22_X1 U1478 ( .A1(n4636), .A2(\REGISTERS[4][17] ), .B1(n4633), .B2(
        \REGISTERS[5][17] ), .ZN(n1980) );
  OAI221_X1 U1479 ( .B1(n1030), .B2(n4690), .C1(n1031), .C2(n4687), .A(n1954), 
        .ZN(n1949) );
  AOI22_X1 U1480 ( .A1(n4684), .A2(\REGISTERS[20][18] ), .B1(n4681), .B2(
        \REGISTERS[21][18] ), .ZN(n1954) );
  OAI221_X1 U1481 ( .B1(n1046), .B2(n4642), .C1(n1047), .C2(n4639), .A(n1962), 
        .ZN(n1957) );
  AOI22_X1 U1482 ( .A1(n4636), .A2(\REGISTERS[4][18] ), .B1(n4633), .B2(
        \REGISTERS[5][18] ), .ZN(n1962) );
  OAI221_X1 U1483 ( .B1(n996), .B2(n4690), .C1(n997), .C2(n4687), .A(n1936), 
        .ZN(n1931) );
  AOI22_X1 U1484 ( .A1(n4684), .A2(\REGISTERS[20][19] ), .B1(n4681), .B2(
        \REGISTERS[21][19] ), .ZN(n1936) );
  OAI221_X1 U1485 ( .B1(n1012), .B2(n4642), .C1(n1013), .C2(n4639), .A(n1944), 
        .ZN(n1939) );
  AOI22_X1 U1486 ( .A1(n4636), .A2(\REGISTERS[4][19] ), .B1(n4633), .B2(
        \REGISTERS[5][19] ), .ZN(n1944) );
  OAI221_X1 U1487 ( .B1(n962), .B2(n4690), .C1(n963), .C2(n4687), .A(n1918), 
        .ZN(n1913) );
  AOI22_X1 U1488 ( .A1(n4684), .A2(\REGISTERS[20][20] ), .B1(n4681), .B2(
        \REGISTERS[21][20] ), .ZN(n1918) );
  OAI221_X1 U1489 ( .B1(n978), .B2(n4642), .C1(n979), .C2(n4639), .A(n1926), 
        .ZN(n1921) );
  AOI22_X1 U1490 ( .A1(n4636), .A2(\REGISTERS[4][20] ), .B1(n4633), .B2(
        \REGISTERS[5][20] ), .ZN(n1926) );
  OAI221_X1 U1491 ( .B1(n928), .B2(n4690), .C1(n929), .C2(n4687), .A(n1900), 
        .ZN(n1895) );
  AOI22_X1 U1492 ( .A1(n4684), .A2(\REGISTERS[20][21] ), .B1(n4681), .B2(
        \REGISTERS[21][21] ), .ZN(n1900) );
  OAI221_X1 U1493 ( .B1(n944), .B2(n4642), .C1(n945), .C2(n4639), .A(n1908), 
        .ZN(n1903) );
  AOI22_X1 U1494 ( .A1(n4636), .A2(\REGISTERS[4][21] ), .B1(n4633), .B2(
        \REGISTERS[5][21] ), .ZN(n1908) );
  OAI221_X1 U1495 ( .B1(n4773), .B2(n1654), .C1(n4770), .C2(n1655), .A(n1656), 
        .ZN(n1632) );
  AOI22_X1 U1496 ( .A1(\REGISTERS[16][0] ), .A2(n4767), .B1(\REGISTERS[17][0] ), .B2(n4764), .ZN(n1656) );
  OAI221_X1 U1497 ( .B1(n4773), .B2(n1611), .C1(n4770), .C2(n1612), .A(n1613), 
        .ZN(n1598) );
  AOI22_X1 U1498 ( .A1(\REGISTERS[16][1] ), .A2(n4767), .B1(\REGISTERS[17][1] ), .B2(n4764), .ZN(n1613) );
  OAI221_X1 U1499 ( .B1(n4773), .B2(n1577), .C1(n4770), .C2(n1578), .A(n1579), 
        .ZN(n1564) );
  AOI22_X1 U1500 ( .A1(\REGISTERS[16][2] ), .A2(n4767), .B1(\REGISTERS[17][2] ), .B2(n4764), .ZN(n1579) );
  OAI221_X1 U1501 ( .B1(n4773), .B2(n1543), .C1(n4770), .C2(n1544), .A(n1545), 
        .ZN(n1530) );
  AOI22_X1 U1502 ( .A1(\REGISTERS[16][3] ), .A2(n4767), .B1(\REGISTERS[17][3] ), .B2(n4764), .ZN(n1545) );
  OAI221_X1 U1503 ( .B1(n4773), .B2(n1509), .C1(n4770), .C2(n1510), .A(n1511), 
        .ZN(n1496) );
  AOI22_X1 U1504 ( .A1(\REGISTERS[16][4] ), .A2(n4767), .B1(\REGISTERS[17][4] ), .B2(n4764), .ZN(n1511) );
  OAI221_X1 U1505 ( .B1(n4773), .B2(n1475), .C1(n4770), .C2(n1476), .A(n1477), 
        .ZN(n1462) );
  AOI22_X1 U1506 ( .A1(\REGISTERS[16][5] ), .A2(n4767), .B1(\REGISTERS[17][5] ), .B2(n4764), .ZN(n1477) );
  OAI221_X1 U1507 ( .B1(n4773), .B2(n1441), .C1(n4770), .C2(n1442), .A(n1443), 
        .ZN(n1428) );
  AOI22_X1 U1508 ( .A1(\REGISTERS[16][6] ), .A2(n4767), .B1(\REGISTERS[17][6] ), .B2(n4764), .ZN(n1443) );
  OAI221_X1 U1509 ( .B1(n4773), .B2(n1407), .C1(n4770), .C2(n1408), .A(n1409), 
        .ZN(n1394) );
  AOI22_X1 U1510 ( .A1(\REGISTERS[16][7] ), .A2(n4767), .B1(\REGISTERS[17][7] ), .B2(n4764), .ZN(n1409) );
  OAI221_X1 U1511 ( .B1(n4773), .B2(n1373), .C1(n4770), .C2(n1374), .A(n1375), 
        .ZN(n1360) );
  AOI22_X1 U1512 ( .A1(\REGISTERS[16][8] ), .A2(n4767), .B1(\REGISTERS[17][8] ), .B2(n4764), .ZN(n1375) );
  OAI221_X1 U1513 ( .B1(n4773), .B2(n1339), .C1(n4770), .C2(n1340), .A(n1341), 
        .ZN(n1326) );
  AOI22_X1 U1514 ( .A1(\REGISTERS[16][9] ), .A2(n4767), .B1(\REGISTERS[17][9] ), .B2(n4764), .ZN(n1341) );
  OAI221_X1 U1515 ( .B1(n4773), .B2(n1305), .C1(n4770), .C2(n1306), .A(n1307), 
        .ZN(n1292) );
  AOI22_X1 U1516 ( .A1(\REGISTERS[16][10] ), .A2(n4767), .B1(
        \REGISTERS[17][10] ), .B2(n4764), .ZN(n1307) );
  OAI221_X1 U1517 ( .B1(n4773), .B2(n1271), .C1(n4771), .C2(n1272), .A(n1273), 
        .ZN(n1258) );
  AOI22_X1 U1518 ( .A1(\REGISTERS[16][11] ), .A2(n4767), .B1(
        \REGISTERS[17][11] ), .B2(n4764), .ZN(n1273) );
  OAI221_X1 U1519 ( .B1(n4774), .B2(n1237), .C1(n4771), .C2(n1238), .A(n1239), 
        .ZN(n1224) );
  AOI22_X1 U1520 ( .A1(\REGISTERS[16][12] ), .A2(n4768), .B1(
        \REGISTERS[17][12] ), .B2(n4765), .ZN(n1239) );
  OAI221_X1 U1521 ( .B1(n4774), .B2(n1203), .C1(n4771), .C2(n1204), .A(n1205), 
        .ZN(n1190) );
  AOI22_X1 U1522 ( .A1(\REGISTERS[16][13] ), .A2(n4768), .B1(
        \REGISTERS[17][13] ), .B2(n4765), .ZN(n1205) );
  OAI221_X1 U1523 ( .B1(n4774), .B2(n1169), .C1(n4771), .C2(n1170), .A(n1171), 
        .ZN(n1156) );
  AOI22_X1 U1524 ( .A1(\REGISTERS[16][14] ), .A2(n4768), .B1(
        \REGISTERS[17][14] ), .B2(n4765), .ZN(n1171) );
  OAI221_X1 U1525 ( .B1(n4774), .B2(n1135), .C1(n4771), .C2(n1136), .A(n1137), 
        .ZN(n1122) );
  AOI22_X1 U1526 ( .A1(\REGISTERS[16][15] ), .A2(n4768), .B1(
        \REGISTERS[17][15] ), .B2(n4765), .ZN(n1137) );
  OAI221_X1 U1527 ( .B1(n4774), .B2(n1101), .C1(n4771), .C2(n1102), .A(n1103), 
        .ZN(n1088) );
  AOI22_X1 U1528 ( .A1(\REGISTERS[16][16] ), .A2(n4768), .B1(
        \REGISTERS[17][16] ), .B2(n4765), .ZN(n1103) );
  OAI221_X1 U1529 ( .B1(n4774), .B2(n1067), .C1(n4771), .C2(n1068), .A(n1069), 
        .ZN(n1054) );
  AOI22_X1 U1530 ( .A1(\REGISTERS[16][17] ), .A2(n4768), .B1(
        \REGISTERS[17][17] ), .B2(n4765), .ZN(n1069) );
  OAI221_X1 U1531 ( .B1(n4774), .B2(n1033), .C1(n4771), .C2(n1034), .A(n1035), 
        .ZN(n1020) );
  AOI22_X1 U1532 ( .A1(\REGISTERS[16][18] ), .A2(n4768), .B1(
        \REGISTERS[17][18] ), .B2(n4765), .ZN(n1035) );
  OAI221_X1 U1533 ( .B1(n4774), .B2(n999), .C1(n4771), .C2(n1000), .A(n1001), 
        .ZN(n986) );
  AOI22_X1 U1534 ( .A1(\REGISTERS[16][19] ), .A2(n4768), .B1(
        \REGISTERS[17][19] ), .B2(n4765), .ZN(n1001) );
  OAI221_X1 U1535 ( .B1(n4774), .B2(n965), .C1(n4771), .C2(n966), .A(n967), 
        .ZN(n952) );
  AOI22_X1 U1536 ( .A1(\REGISTERS[16][20] ), .A2(n4768), .B1(
        \REGISTERS[17][20] ), .B2(n4765), .ZN(n967) );
  OAI221_X1 U1537 ( .B1(n4774), .B2(n931), .C1(n4771), .C2(n932), .A(n933), 
        .ZN(n918) );
  AOI22_X1 U1538 ( .A1(\REGISTERS[16][21] ), .A2(n4768), .B1(
        \REGISTERS[17][21] ), .B2(n4765), .ZN(n933) );
  OAI221_X1 U1539 ( .B1(n4774), .B2(n897), .C1(n4772), .C2(n898), .A(n899), 
        .ZN(n884) );
  AOI22_X1 U1540 ( .A1(\REGISTERS[16][22] ), .A2(n4768), .B1(
        \REGISTERS[17][22] ), .B2(n4765), .ZN(n899) );
  OAI221_X1 U1541 ( .B1(n4774), .B2(n863), .C1(n4772), .C2(n864), .A(n865), 
        .ZN(n850) );
  AOI22_X1 U1542 ( .A1(\REGISTERS[16][23] ), .A2(n4768), .B1(
        \REGISTERS[17][23] ), .B2(n4765), .ZN(n865) );
  OAI221_X1 U1543 ( .B1(n1271), .B2(n4678), .C1(n1272), .C2(n4675), .A(n2081), 
        .ZN(n2074) );
  AOI22_X1 U1544 ( .A1(n4672), .A2(\REGISTERS[16][11] ), .B1(n4669), .B2(
        \REGISTERS[17][11] ), .ZN(n2081) );
  OAI221_X1 U1545 ( .B1(n1237), .B2(n4678), .C1(n1238), .C2(n4675), .A(n2063), 
        .ZN(n2056) );
  AOI22_X1 U1546 ( .A1(n4672), .A2(\REGISTERS[16][12] ), .B1(n4669), .B2(
        \REGISTERS[17][12] ), .ZN(n2063) );
  OAI221_X1 U1547 ( .B1(n1203), .B2(n4678), .C1(n1204), .C2(n4675), .A(n2045), 
        .ZN(n2038) );
  AOI22_X1 U1548 ( .A1(n4672), .A2(\REGISTERS[16][13] ), .B1(n4669), .B2(
        \REGISTERS[17][13] ), .ZN(n2045) );
  OAI221_X1 U1549 ( .B1(n1169), .B2(n4678), .C1(n1170), .C2(n4675), .A(n2027), 
        .ZN(n2020) );
  AOI22_X1 U1550 ( .A1(n4672), .A2(\REGISTERS[16][14] ), .B1(n4669), .B2(
        \REGISTERS[17][14] ), .ZN(n2027) );
  OAI221_X1 U1551 ( .B1(n1135), .B2(n4678), .C1(n1136), .C2(n4675), .A(n2009), 
        .ZN(n2002) );
  AOI22_X1 U1552 ( .A1(n4672), .A2(\REGISTERS[16][15] ), .B1(n4669), .B2(
        \REGISTERS[17][15] ), .ZN(n2009) );
  OAI221_X1 U1553 ( .B1(n1101), .B2(n4678), .C1(n1102), .C2(n4675), .A(n1991), 
        .ZN(n1984) );
  AOI22_X1 U1554 ( .A1(n4672), .A2(\REGISTERS[16][16] ), .B1(n4669), .B2(
        \REGISTERS[17][16] ), .ZN(n1991) );
  OAI221_X1 U1555 ( .B1(n1067), .B2(n4678), .C1(n1068), .C2(n4675), .A(n1973), 
        .ZN(n1966) );
  AOI22_X1 U1556 ( .A1(n4672), .A2(\REGISTERS[16][17] ), .B1(n4669), .B2(
        \REGISTERS[17][17] ), .ZN(n1973) );
  OAI221_X1 U1557 ( .B1(n1033), .B2(n4678), .C1(n1034), .C2(n4675), .A(n1955), 
        .ZN(n1948) );
  AOI22_X1 U1558 ( .A1(n4672), .A2(\REGISTERS[16][18] ), .B1(n4669), .B2(
        \REGISTERS[17][18] ), .ZN(n1955) );
  OAI221_X1 U1559 ( .B1(n999), .B2(n4678), .C1(n1000), .C2(n4675), .A(n1937), 
        .ZN(n1930) );
  AOI22_X1 U1560 ( .A1(n4672), .A2(\REGISTERS[16][19] ), .B1(n4669), .B2(
        \REGISTERS[17][19] ), .ZN(n1937) );
  OAI221_X1 U1561 ( .B1(n965), .B2(n4678), .C1(n966), .C2(n4675), .A(n1919), 
        .ZN(n1912) );
  AOI22_X1 U1562 ( .A1(n4672), .A2(\REGISTERS[16][20] ), .B1(n4669), .B2(
        \REGISTERS[17][20] ), .ZN(n1919) );
  OAI221_X1 U1563 ( .B1(n931), .B2(n4678), .C1(n932), .C2(n4675), .A(n1901), 
        .ZN(n1894) );
  AOI22_X1 U1564 ( .A1(n4672), .A2(\REGISTERS[16][21] ), .B1(n4669), .B2(
        \REGISTERS[17][21] ), .ZN(n1901) );
  NAND2_X1 U1565 ( .A1(n5080), .A2(ENABLE), .ZN(n525) );
  AND3_X1 U1566 ( .A1(n1675), .A2(n1676), .A3(ADD_RD2[2]), .ZN(n1640) );
  AND3_X1 U1567 ( .A1(n1675), .A2(n2301), .A3(ADD_RD1[2]), .ZN(n2278) );
  AOI22_X1 U1568 ( .A1(\REGISTERS[0][24] ), .A2(n4721), .B1(\REGISTERS[1][24] ), .B2(n4718), .ZN(n847) );
  AOI22_X1 U1569 ( .A1(\REGISTERS[0][25] ), .A2(n4721), .B1(\REGISTERS[1][25] ), .B2(n4718), .ZN(n813) );
  AOI22_X1 U1570 ( .A1(\REGISTERS[0][26] ), .A2(n4721), .B1(\REGISTERS[1][26] ), .B2(n4718), .ZN(n779) );
  AOI22_X1 U1571 ( .A1(\REGISTERS[0][27] ), .A2(n4721), .B1(\REGISTERS[1][27] ), .B2(n4718), .ZN(n745) );
  AOI22_X1 U1572 ( .A1(\REGISTERS[0][28] ), .A2(n4721), .B1(\REGISTERS[1][28] ), .B2(n4718), .ZN(n711) );
  AOI22_X1 U1573 ( .A1(\REGISTERS[0][29] ), .A2(n4721), .B1(\REGISTERS[1][29] ), .B2(n4718), .ZN(n677) );
  AOI22_X1 U1574 ( .A1(\REGISTERS[0][30] ), .A2(n4721), .B1(\REGISTERS[1][30] ), .B2(n4718), .ZN(n643) );
  AOI22_X1 U1575 ( .A1(\REGISTERS[0][31] ), .A2(n4721), .B1(\REGISTERS[1][31] ), .B2(n4718), .ZN(n607) );
  AOI22_X1 U1576 ( .A1(\REGISTERS[0][0] ), .A2(n4719), .B1(\REGISTERS[1][0] ), 
        .B2(n4716), .ZN(n1679) );
  AOI22_X1 U1577 ( .A1(\REGISTERS[0][1] ), .A2(n4719), .B1(\REGISTERS[1][1] ), 
        .B2(n4716), .ZN(n1629) );
  AOI22_X1 U1578 ( .A1(\REGISTERS[0][2] ), .A2(n4719), .B1(\REGISTERS[1][2] ), 
        .B2(n4716), .ZN(n1595) );
  AOI22_X1 U1579 ( .A1(\REGISTERS[0][3] ), .A2(n4719), .B1(\REGISTERS[1][3] ), 
        .B2(n4716), .ZN(n1561) );
  AOI22_X1 U1580 ( .A1(\REGISTERS[0][4] ), .A2(n4719), .B1(\REGISTERS[1][4] ), 
        .B2(n4716), .ZN(n1527) );
  AOI22_X1 U1581 ( .A1(\REGISTERS[0][5] ), .A2(n4719), .B1(\REGISTERS[1][5] ), 
        .B2(n4716), .ZN(n1493) );
  AOI22_X1 U1582 ( .A1(\REGISTERS[0][6] ), .A2(n4719), .B1(\REGISTERS[1][6] ), 
        .B2(n4716), .ZN(n1459) );
  AOI22_X1 U1583 ( .A1(\REGISTERS[0][7] ), .A2(n4719), .B1(\REGISTERS[1][7] ), 
        .B2(n4716), .ZN(n1425) );
  AOI22_X1 U1584 ( .A1(\REGISTERS[0][8] ), .A2(n4719), .B1(\REGISTERS[1][8] ), 
        .B2(n4716), .ZN(n1391) );
  AOI22_X1 U1585 ( .A1(\REGISTERS[0][9] ), .A2(n4719), .B1(\REGISTERS[1][9] ), 
        .B2(n4716), .ZN(n1357) );
  AOI22_X1 U1586 ( .A1(\REGISTERS[0][10] ), .A2(n4719), .B1(\REGISTERS[1][10] ), .B2(n4716), .ZN(n1323) );
  AOI22_X1 U1587 ( .A1(\REGISTERS[0][11] ), .A2(n4719), .B1(\REGISTERS[1][11] ), .B2(n4716), .ZN(n1289) );
  AOI22_X1 U1588 ( .A1(\REGISTERS[0][12] ), .A2(n4720), .B1(\REGISTERS[1][12] ), .B2(n4717), .ZN(n1255) );
  AOI22_X1 U1589 ( .A1(\REGISTERS[0][13] ), .A2(n4720), .B1(\REGISTERS[1][13] ), .B2(n4717), .ZN(n1221) );
  AOI22_X1 U1590 ( .A1(\REGISTERS[0][14] ), .A2(n4720), .B1(\REGISTERS[1][14] ), .B2(n4717), .ZN(n1187) );
  AOI22_X1 U1591 ( .A1(\REGISTERS[0][15] ), .A2(n4720), .B1(\REGISTERS[1][15] ), .B2(n4717), .ZN(n1153) );
  AOI22_X1 U1592 ( .A1(\REGISTERS[0][16] ), .A2(n4720), .B1(\REGISTERS[1][16] ), .B2(n4717), .ZN(n1119) );
  AOI22_X1 U1593 ( .A1(\REGISTERS[0][17] ), .A2(n4720), .B1(\REGISTERS[1][17] ), .B2(n4717), .ZN(n1085) );
  AOI22_X1 U1594 ( .A1(\REGISTERS[0][18] ), .A2(n4720), .B1(\REGISTERS[1][18] ), .B2(n4717), .ZN(n1051) );
  AOI22_X1 U1595 ( .A1(\REGISTERS[0][19] ), .A2(n4720), .B1(\REGISTERS[1][19] ), .B2(n4717), .ZN(n1017) );
  AOI22_X1 U1596 ( .A1(\REGISTERS[0][20] ), .A2(n4720), .B1(\REGISTERS[1][20] ), .B2(n4717), .ZN(n983) );
  AOI22_X1 U1597 ( .A1(\REGISTERS[0][21] ), .A2(n4720), .B1(\REGISTERS[1][21] ), .B2(n4717), .ZN(n949) );
  AOI22_X1 U1598 ( .A1(\REGISTERS[0][22] ), .A2(n4720), .B1(\REGISTERS[1][22] ), .B2(n4717), .ZN(n915) );
  AOI22_X1 U1599 ( .A1(\REGISTERS[0][23] ), .A2(n4720), .B1(\REGISTERS[1][23] ), .B2(n4717), .ZN(n881) );
  AOI22_X1 U1600 ( .A1(n4623), .A2(\REGISTERS[0][0] ), .B1(n4620), .B2(
        \REGISTERS[1][0] ), .ZN(n2302) );
  AOI22_X1 U1601 ( .A1(n4623), .A2(\REGISTERS[0][1] ), .B1(n4620), .B2(
        \REGISTERS[1][1] ), .ZN(n2269) );
  AOI22_X1 U1602 ( .A1(n4623), .A2(\REGISTERS[0][2] ), .B1(n4620), .B2(
        \REGISTERS[1][2] ), .ZN(n2251) );
  AOI22_X1 U1603 ( .A1(n4623), .A2(\REGISTERS[0][3] ), .B1(n4620), .B2(
        \REGISTERS[1][3] ), .ZN(n2233) );
  AOI22_X1 U1604 ( .A1(n4623), .A2(\REGISTERS[0][4] ), .B1(n4620), .B2(
        \REGISTERS[1][4] ), .ZN(n2215) );
  AOI22_X1 U1605 ( .A1(n4623), .A2(\REGISTERS[0][5] ), .B1(n4620), .B2(
        \REGISTERS[1][5] ), .ZN(n2197) );
  AOI22_X1 U1606 ( .A1(n4623), .A2(\REGISTERS[0][6] ), .B1(n4620), .B2(
        \REGISTERS[1][6] ), .ZN(n2179) );
  AOI22_X1 U1607 ( .A1(n4623), .A2(\REGISTERS[0][7] ), .B1(n4620), .B2(
        \REGISTERS[1][7] ), .ZN(n2161) );
  AOI22_X1 U1608 ( .A1(n4623), .A2(\REGISTERS[0][8] ), .B1(n4620), .B2(
        \REGISTERS[1][8] ), .ZN(n2143) );
  AOI22_X1 U1609 ( .A1(n4623), .A2(\REGISTERS[0][9] ), .B1(n4620), .B2(
        \REGISTERS[1][9] ), .ZN(n2125) );
  AOI22_X1 U1610 ( .A1(n4623), .A2(\REGISTERS[0][10] ), .B1(n4620), .B2(
        \REGISTERS[1][10] ), .ZN(n2107) );
  AOI22_X1 U1611 ( .A1(n4624), .A2(\REGISTERS[0][11] ), .B1(n4621), .B2(
        \REGISTERS[1][11] ), .ZN(n2089) );
  AOI22_X1 U1612 ( .A1(n4624), .A2(\REGISTERS[0][12] ), .B1(n4621), .B2(
        \REGISTERS[1][12] ), .ZN(n2071) );
  AOI22_X1 U1613 ( .A1(n4624), .A2(\REGISTERS[0][13] ), .B1(n4621), .B2(
        \REGISTERS[1][13] ), .ZN(n2053) );
  AOI22_X1 U1614 ( .A1(n4624), .A2(\REGISTERS[0][14] ), .B1(n4621), .B2(
        \REGISTERS[1][14] ), .ZN(n2035) );
  AOI22_X1 U1615 ( .A1(n4624), .A2(\REGISTERS[0][15] ), .B1(n4621), .B2(
        \REGISTERS[1][15] ), .ZN(n2017) );
  AOI22_X1 U1616 ( .A1(n4624), .A2(\REGISTERS[0][16] ), .B1(n4621), .B2(
        \REGISTERS[1][16] ), .ZN(n1999) );
  AOI22_X1 U1617 ( .A1(n4624), .A2(\REGISTERS[0][17] ), .B1(n4621), .B2(
        \REGISTERS[1][17] ), .ZN(n1981) );
  AOI22_X1 U1618 ( .A1(n4624), .A2(\REGISTERS[0][18] ), .B1(n4621), .B2(
        \REGISTERS[1][18] ), .ZN(n1963) );
  AOI22_X1 U1619 ( .A1(n4624), .A2(\REGISTERS[0][19] ), .B1(n4621), .B2(
        \REGISTERS[1][19] ), .ZN(n1945) );
  AOI22_X1 U1620 ( .A1(n4624), .A2(\REGISTERS[0][20] ), .B1(n4621), .B2(
        \REGISTERS[1][20] ), .ZN(n1927) );
  AOI22_X1 U1621 ( .A1(n4624), .A2(\REGISTERS[0][21] ), .B1(n4621), .B2(
        \REGISTERS[1][21] ), .ZN(n1909) );
  AOI22_X1 U1622 ( .A1(n4625), .A2(\REGISTERS[0][22] ), .B1(n4622), .B2(
        \REGISTERS[1][22] ), .ZN(n1891) );
  AOI22_X1 U1623 ( .A1(n4625), .A2(\REGISTERS[0][23] ), .B1(n4622), .B2(
        \REGISTERS[1][23] ), .ZN(n1873) );
  AOI22_X1 U1624 ( .A1(n4625), .A2(\REGISTERS[0][24] ), .B1(n4622), .B2(
        \REGISTERS[1][24] ), .ZN(n1855) );
  AOI22_X1 U1625 ( .A1(n4625), .A2(\REGISTERS[0][25] ), .B1(n4622), .B2(
        \REGISTERS[1][25] ), .ZN(n1837) );
  AOI22_X1 U1626 ( .A1(n4625), .A2(\REGISTERS[0][26] ), .B1(n4622), .B2(
        \REGISTERS[1][26] ), .ZN(n1819) );
  AOI22_X1 U1627 ( .A1(n4625), .A2(\REGISTERS[0][27] ), .B1(n4622), .B2(
        \REGISTERS[1][27] ), .ZN(n1801) );
  AOI22_X1 U1628 ( .A1(n4625), .A2(\REGISTERS[0][28] ), .B1(n4622), .B2(
        \REGISTERS[1][28] ), .ZN(n1783) );
  AOI22_X1 U1629 ( .A1(n4625), .A2(\REGISTERS[0][29] ), .B1(n4622), .B2(
        \REGISTERS[1][29] ), .ZN(n1765) );
  AOI22_X1 U1630 ( .A1(n4625), .A2(\REGISTERS[0][30] ), .B1(n4622), .B2(
        \REGISTERS[1][30] ), .ZN(n1747) );
  AOI22_X1 U1631 ( .A1(n4625), .A2(\REGISTERS[0][31] ), .B1(n4622), .B2(
        \REGISTERS[1][31] ), .ZN(n1727) );
  AND3_X1 U1632 ( .A1(ADD_RD2[4]), .A2(n1657), .A3(ADD_RD2[0]), .ZN(n1652) );
  AND3_X1 U1633 ( .A1(ADD_RD1[4]), .A2(n2289), .A3(ADD_RD1[0]), .ZN(n2286) );
  AND3_X1 U1634 ( .A1(n1648), .A2(n1657), .A3(ADD_RD2[4]), .ZN(n1653) );
  AND3_X1 U1635 ( .A1(n2284), .A2(n2289), .A3(ADD_RD1[4]), .ZN(n2287) );
  OR2_X1 U1636 ( .A1(RD2), .A2(n525), .ZN(n4608) );
  OR2_X1 U1637 ( .A1(RD1), .A2(n525), .ZN(n4612) );
  AND3_X1 U1638 ( .A1(ADD_RD2[4]), .A2(n1648), .A3(ADD_RD2[3]), .ZN(n1641) );
  AND3_X1 U1639 ( .A1(ADD_RD1[4]), .A2(n2284), .A3(ADD_RD1[3]), .ZN(n2279) );
  AND3_X1 U1640 ( .A1(ADD_RD2[0]), .A2(ADD_RD2[4]), .A3(ADD_RD2[3]), .ZN(n1639) );
  AND3_X1 U1641 ( .A1(ADD_RD1[0]), .A2(ADD_RD1[4]), .A3(ADD_RD1[3]), .ZN(n2277) );
  INV_X1 U1642 ( .A(ADD_RD2[3]), .ZN(n1657) );
  INV_X1 U1643 ( .A(ADD_RD2[0]), .ZN(n1648) );
  INV_X1 U1644 ( .A(ADD_RD1[3]), .ZN(n2289) );
  INV_X1 U1645 ( .A(ADD_RD1[0]), .ZN(n2284) );
  AND2_X1 U1646 ( .A1(WR), .A2(ENABLE), .ZN(n535) );
  AND2_X1 U1647 ( .A1(DATAIN[31]), .A2(n5080), .ZN(n4352) );
  AND2_X1 U1648 ( .A1(DATAIN[0]), .A2(n5081), .ZN(n4480) );
  AND2_X1 U1649 ( .A1(DATAIN[1]), .A2(n5081), .ZN(n4476) );
  AND2_X1 U1650 ( .A1(DATAIN[2]), .A2(n5081), .ZN(n4472) );
  AND2_X1 U1651 ( .A1(DATAIN[3]), .A2(n5081), .ZN(n4468) );
  AND2_X1 U1652 ( .A1(DATAIN[4]), .A2(n5081), .ZN(n4464) );
  AND2_X1 U1653 ( .A1(DATAIN[5]), .A2(n5081), .ZN(n4460) );
  AND2_X1 U1654 ( .A1(DATAIN[6]), .A2(n5081), .ZN(n4456) );
  AND2_X1 U1655 ( .A1(DATAIN[7]), .A2(n5081), .ZN(n4452) );
  AND2_X1 U1656 ( .A1(DATAIN[8]), .A2(n5081), .ZN(n4448) );
  AND2_X1 U1657 ( .A1(DATAIN[9]), .A2(n5081), .ZN(n4444) );
  AND2_X1 U1658 ( .A1(DATAIN[10]), .A2(n5081), .ZN(n4440) );
  AND2_X1 U1659 ( .A1(DATAIN[11]), .A2(n5081), .ZN(n4436) );
  AND2_X1 U1660 ( .A1(DATAIN[12]), .A2(n5081), .ZN(n4432) );
  AND2_X1 U1661 ( .A1(DATAIN[13]), .A2(n5081), .ZN(n4428) );
  AND2_X1 U1662 ( .A1(DATAIN[14]), .A2(n5081), .ZN(n4424) );
  AND2_X1 U1663 ( .A1(DATAIN[15]), .A2(n5081), .ZN(n4420) );
  AND2_X1 U1664 ( .A1(DATAIN[16]), .A2(n5081), .ZN(n4416) );
  AND2_X1 U1665 ( .A1(DATAIN[17]), .A2(n5081), .ZN(n4412) );
  AND2_X1 U1666 ( .A1(DATAIN[18]), .A2(n5082), .ZN(n4408) );
  AND2_X1 U1667 ( .A1(DATAIN[19]), .A2(n5082), .ZN(n4404) );
  AND2_X1 U1668 ( .A1(DATAIN[20]), .A2(n5082), .ZN(n4400) );
  AND2_X1 U1669 ( .A1(DATAIN[21]), .A2(n5082), .ZN(n4396) );
  AND2_X1 U1670 ( .A1(DATAIN[22]), .A2(n5082), .ZN(n4392) );
  AND2_X1 U1671 ( .A1(DATAIN[23]), .A2(n5082), .ZN(n4388) );
  AND2_X1 U1672 ( .A1(DATAIN[24]), .A2(n5082), .ZN(n4384) );
  AND2_X1 U1673 ( .A1(DATAIN[25]), .A2(n5082), .ZN(n4380) );
  AND2_X1 U1674 ( .A1(DATAIN[26]), .A2(n5082), .ZN(n4376) );
  AND2_X1 U1675 ( .A1(DATAIN[27]), .A2(n5082), .ZN(n4372) );
  AND2_X1 U1676 ( .A1(DATAIN[28]), .A2(n5082), .ZN(n4368) );
  AND2_X1 U1677 ( .A1(DATAIN[29]), .A2(n5082), .ZN(n4364) );
  AND2_X1 U1678 ( .A1(DATAIN[30]), .A2(n5082), .ZN(n4360) );
  INV_X1 U1679 ( .A(ADD_RD2[1]), .ZN(n1676) );
  INV_X1 U1680 ( .A(\REGISTERS[30][0] ), .ZN(n1636) );
  INV_X1 U1681 ( .A(\REGISTERS[26][0] ), .ZN(n1643) );
  INV_X1 U1682 ( .A(\REGISTERS[22][0] ), .ZN(n1649) );
  INV_X1 U1683 ( .A(\REGISTERS[18][0] ), .ZN(n1654) );
  INV_X1 U1684 ( .A(\REGISTERS[14][0] ), .ZN(n1662) );
  INV_X1 U1685 ( .A(\REGISTERS[10][0] ), .ZN(n1667) );
  INV_X1 U1686 ( .A(\REGISTERS[6][0] ), .ZN(n1670) );
  INV_X1 U1687 ( .A(\REGISTERS[2][0] ), .ZN(n1677) );
  INV_X1 U1688 ( .A(\REGISTERS[30][1] ), .ZN(n1602) );
  INV_X1 U1689 ( .A(\REGISTERS[26][1] ), .ZN(n1605) );
  INV_X1 U1690 ( .A(\REGISTERS[22][1] ), .ZN(n1608) );
  INV_X1 U1691 ( .A(\REGISTERS[18][1] ), .ZN(n1611) );
  INV_X1 U1692 ( .A(\REGISTERS[14][1] ), .ZN(n1618) );
  INV_X1 U1693 ( .A(\REGISTERS[10][1] ), .ZN(n1621) );
  INV_X1 U1694 ( .A(\REGISTERS[6][1] ), .ZN(n1624) );
  INV_X1 U1695 ( .A(\REGISTERS[2][1] ), .ZN(n1627) );
  INV_X1 U1696 ( .A(\REGISTERS[30][2] ), .ZN(n1568) );
  INV_X1 U1697 ( .A(\REGISTERS[26][2] ), .ZN(n1571) );
  INV_X1 U1698 ( .A(\REGISTERS[22][2] ), .ZN(n1574) );
  INV_X1 U1699 ( .A(\REGISTERS[18][2] ), .ZN(n1577) );
  INV_X1 U1700 ( .A(\REGISTERS[14][2] ), .ZN(n1584) );
  INV_X1 U1701 ( .A(\REGISTERS[10][2] ), .ZN(n1587) );
  INV_X1 U1702 ( .A(\REGISTERS[6][2] ), .ZN(n1590) );
  INV_X1 U1703 ( .A(\REGISTERS[2][2] ), .ZN(n1593) );
  INV_X1 U1704 ( .A(\REGISTERS[30][3] ), .ZN(n1534) );
  INV_X1 U1705 ( .A(\REGISTERS[26][3] ), .ZN(n1537) );
  INV_X1 U1706 ( .A(\REGISTERS[22][3] ), .ZN(n1540) );
  INV_X1 U1707 ( .A(\REGISTERS[18][3] ), .ZN(n1543) );
  INV_X1 U1708 ( .A(\REGISTERS[14][3] ), .ZN(n1550) );
  INV_X1 U1709 ( .A(\REGISTERS[10][3] ), .ZN(n1553) );
  INV_X1 U1710 ( .A(\REGISTERS[6][3] ), .ZN(n1556) );
  INV_X1 U1711 ( .A(\REGISTERS[2][3] ), .ZN(n1559) );
  INV_X1 U1712 ( .A(\REGISTERS[30][4] ), .ZN(n1500) );
  INV_X1 U1713 ( .A(\REGISTERS[26][4] ), .ZN(n1503) );
  INV_X1 U1714 ( .A(\REGISTERS[22][4] ), .ZN(n1506) );
  INV_X1 U1715 ( .A(\REGISTERS[18][4] ), .ZN(n1509) );
  INV_X1 U1716 ( .A(\REGISTERS[14][4] ), .ZN(n1516) );
  INV_X1 U1717 ( .A(\REGISTERS[10][4] ), .ZN(n1519) );
  INV_X1 U1718 ( .A(\REGISTERS[6][4] ), .ZN(n1522) );
  INV_X1 U1719 ( .A(\REGISTERS[2][4] ), .ZN(n1525) );
  INV_X1 U1720 ( .A(\REGISTERS[30][5] ), .ZN(n1466) );
  INV_X1 U1721 ( .A(\REGISTERS[26][5] ), .ZN(n1469) );
  INV_X1 U1722 ( .A(\REGISTERS[22][5] ), .ZN(n1472) );
  INV_X1 U1723 ( .A(\REGISTERS[18][5] ), .ZN(n1475) );
  INV_X1 U1724 ( .A(\REGISTERS[14][5] ), .ZN(n1482) );
  INV_X1 U1725 ( .A(\REGISTERS[10][5] ), .ZN(n1485) );
  INV_X1 U1726 ( .A(\REGISTERS[6][5] ), .ZN(n1488) );
  INV_X1 U1727 ( .A(\REGISTERS[2][5] ), .ZN(n1491) );
  INV_X1 U1728 ( .A(\REGISTERS[30][6] ), .ZN(n1432) );
  INV_X1 U1729 ( .A(\REGISTERS[26][6] ), .ZN(n1435) );
  INV_X1 U1730 ( .A(\REGISTERS[22][6] ), .ZN(n1438) );
  INV_X1 U1731 ( .A(\REGISTERS[18][6] ), .ZN(n1441) );
  INV_X1 U1732 ( .A(\REGISTERS[14][6] ), .ZN(n1448) );
  INV_X1 U1733 ( .A(\REGISTERS[10][6] ), .ZN(n1451) );
  INV_X1 U1734 ( .A(\REGISTERS[6][6] ), .ZN(n1454) );
  INV_X1 U1735 ( .A(\REGISTERS[2][6] ), .ZN(n1457) );
  INV_X1 U1736 ( .A(\REGISTERS[30][7] ), .ZN(n1398) );
  INV_X1 U1737 ( .A(\REGISTERS[26][7] ), .ZN(n1401) );
  INV_X1 U1738 ( .A(\REGISTERS[22][7] ), .ZN(n1404) );
  INV_X1 U1739 ( .A(\REGISTERS[18][7] ), .ZN(n1407) );
  INV_X1 U1740 ( .A(\REGISTERS[14][7] ), .ZN(n1414) );
  INV_X1 U1741 ( .A(\REGISTERS[10][7] ), .ZN(n1417) );
  INV_X1 U1742 ( .A(\REGISTERS[6][7] ), .ZN(n1420) );
  INV_X1 U1743 ( .A(\REGISTERS[2][7] ), .ZN(n1423) );
  INV_X1 U1744 ( .A(\REGISTERS[30][8] ), .ZN(n1364) );
  INV_X1 U1745 ( .A(\REGISTERS[26][8] ), .ZN(n1367) );
  INV_X1 U1746 ( .A(\REGISTERS[22][8] ), .ZN(n1370) );
  INV_X1 U1747 ( .A(\REGISTERS[18][8] ), .ZN(n1373) );
  INV_X1 U1748 ( .A(\REGISTERS[14][8] ), .ZN(n1380) );
  INV_X1 U1749 ( .A(\REGISTERS[10][8] ), .ZN(n1383) );
  INV_X1 U1750 ( .A(\REGISTERS[6][8] ), .ZN(n1386) );
  INV_X1 U1751 ( .A(\REGISTERS[2][8] ), .ZN(n1389) );
  INV_X1 U1752 ( .A(\REGISTERS[30][9] ), .ZN(n1330) );
  INV_X1 U1753 ( .A(\REGISTERS[26][9] ), .ZN(n1333) );
  INV_X1 U1754 ( .A(\REGISTERS[22][9] ), .ZN(n1336) );
  INV_X1 U1755 ( .A(\REGISTERS[18][9] ), .ZN(n1339) );
  INV_X1 U1756 ( .A(\REGISTERS[14][9] ), .ZN(n1346) );
  INV_X1 U1757 ( .A(\REGISTERS[10][9] ), .ZN(n1349) );
  INV_X1 U1758 ( .A(\REGISTERS[6][9] ), .ZN(n1352) );
  INV_X1 U1759 ( .A(\REGISTERS[2][9] ), .ZN(n1355) );
  INV_X1 U1760 ( .A(\REGISTERS[30][10] ), .ZN(n1296) );
  INV_X1 U1761 ( .A(\REGISTERS[26][10] ), .ZN(n1299) );
  INV_X1 U1762 ( .A(\REGISTERS[22][10] ), .ZN(n1302) );
  INV_X1 U1763 ( .A(\REGISTERS[18][10] ), .ZN(n1305) );
  INV_X1 U1764 ( .A(\REGISTERS[14][10] ), .ZN(n1312) );
  INV_X1 U1765 ( .A(\REGISTERS[10][10] ), .ZN(n1315) );
  INV_X1 U1766 ( .A(\REGISTERS[6][10] ), .ZN(n1318) );
  INV_X1 U1767 ( .A(\REGISTERS[2][10] ), .ZN(n1321) );
  INV_X1 U1768 ( .A(\REGISTERS[30][11] ), .ZN(n1262) );
  INV_X1 U1769 ( .A(\REGISTERS[26][11] ), .ZN(n1265) );
  INV_X1 U1770 ( .A(\REGISTERS[22][11] ), .ZN(n1268) );
  INV_X1 U1771 ( .A(\REGISTERS[18][11] ), .ZN(n1271) );
  INV_X1 U1772 ( .A(\REGISTERS[14][11] ), .ZN(n1278) );
  INV_X1 U1773 ( .A(\REGISTERS[10][11] ), .ZN(n1281) );
  INV_X1 U1774 ( .A(\REGISTERS[6][11] ), .ZN(n1284) );
  INV_X1 U1775 ( .A(\REGISTERS[2][11] ), .ZN(n1287) );
  INV_X1 U1776 ( .A(\REGISTERS[30][12] ), .ZN(n1228) );
  INV_X1 U1777 ( .A(\REGISTERS[26][12] ), .ZN(n1231) );
  INV_X1 U1778 ( .A(\REGISTERS[22][12] ), .ZN(n1234) );
  INV_X1 U1779 ( .A(\REGISTERS[18][12] ), .ZN(n1237) );
  INV_X1 U1780 ( .A(\REGISTERS[14][12] ), .ZN(n1244) );
  INV_X1 U1781 ( .A(\REGISTERS[10][12] ), .ZN(n1247) );
  INV_X1 U1782 ( .A(\REGISTERS[6][12] ), .ZN(n1250) );
  INV_X1 U1783 ( .A(\REGISTERS[2][12] ), .ZN(n1253) );
  INV_X1 U1784 ( .A(\REGISTERS[30][13] ), .ZN(n1194) );
  INV_X1 U1785 ( .A(\REGISTERS[26][13] ), .ZN(n1197) );
  INV_X1 U1786 ( .A(\REGISTERS[22][13] ), .ZN(n1200) );
  INV_X1 U1787 ( .A(\REGISTERS[18][13] ), .ZN(n1203) );
  INV_X1 U1788 ( .A(\REGISTERS[14][13] ), .ZN(n1210) );
  INV_X1 U1789 ( .A(\REGISTERS[10][13] ), .ZN(n1213) );
  INV_X1 U1790 ( .A(\REGISTERS[6][13] ), .ZN(n1216) );
  INV_X1 U1791 ( .A(\REGISTERS[2][13] ), .ZN(n1219) );
  INV_X1 U1792 ( .A(\REGISTERS[30][14] ), .ZN(n1160) );
  INV_X1 U1793 ( .A(\REGISTERS[26][14] ), .ZN(n1163) );
  INV_X1 U1794 ( .A(\REGISTERS[22][14] ), .ZN(n1166) );
  INV_X1 U1795 ( .A(\REGISTERS[18][14] ), .ZN(n1169) );
  INV_X1 U1796 ( .A(\REGISTERS[14][14] ), .ZN(n1176) );
  INV_X1 U1797 ( .A(\REGISTERS[10][14] ), .ZN(n1179) );
  INV_X1 U1798 ( .A(\REGISTERS[6][14] ), .ZN(n1182) );
  INV_X1 U1799 ( .A(\REGISTERS[2][14] ), .ZN(n1185) );
  INV_X1 U1800 ( .A(\REGISTERS[30][15] ), .ZN(n1126) );
  INV_X1 U1801 ( .A(\REGISTERS[26][15] ), .ZN(n1129) );
  INV_X1 U1802 ( .A(\REGISTERS[22][15] ), .ZN(n1132) );
  INV_X1 U1803 ( .A(\REGISTERS[18][15] ), .ZN(n1135) );
  INV_X1 U1804 ( .A(\REGISTERS[14][15] ), .ZN(n1142) );
  INV_X1 U1805 ( .A(\REGISTERS[10][15] ), .ZN(n1145) );
  INV_X1 U1806 ( .A(\REGISTERS[6][15] ), .ZN(n1148) );
  INV_X1 U1807 ( .A(\REGISTERS[2][15] ), .ZN(n1151) );
  INV_X1 U1808 ( .A(\REGISTERS[30][16] ), .ZN(n1092) );
  INV_X1 U1809 ( .A(\REGISTERS[26][16] ), .ZN(n1095) );
  INV_X1 U1810 ( .A(\REGISTERS[22][16] ), .ZN(n1098) );
  INV_X1 U1811 ( .A(\REGISTERS[18][16] ), .ZN(n1101) );
  INV_X1 U1812 ( .A(\REGISTERS[14][16] ), .ZN(n1108) );
  INV_X1 U1813 ( .A(\REGISTERS[10][16] ), .ZN(n1111) );
  INV_X1 U1814 ( .A(\REGISTERS[6][16] ), .ZN(n1114) );
  INV_X1 U1815 ( .A(\REGISTERS[2][16] ), .ZN(n1117) );
  INV_X1 U1816 ( .A(\REGISTERS[30][17] ), .ZN(n1058) );
  INV_X1 U1817 ( .A(\REGISTERS[26][17] ), .ZN(n1061) );
  INV_X1 U1818 ( .A(\REGISTERS[22][17] ), .ZN(n1064) );
  INV_X1 U1819 ( .A(\REGISTERS[18][17] ), .ZN(n1067) );
  INV_X1 U1820 ( .A(\REGISTERS[14][17] ), .ZN(n1074) );
  INV_X1 U1821 ( .A(\REGISTERS[10][17] ), .ZN(n1077) );
  INV_X1 U1822 ( .A(\REGISTERS[6][17] ), .ZN(n1080) );
  INV_X1 U1823 ( .A(\REGISTERS[2][17] ), .ZN(n1083) );
  INV_X1 U1824 ( .A(\REGISTERS[30][18] ), .ZN(n1024) );
  INV_X1 U1825 ( .A(\REGISTERS[26][18] ), .ZN(n1027) );
  INV_X1 U1826 ( .A(\REGISTERS[22][18] ), .ZN(n1030) );
  INV_X1 U1827 ( .A(\REGISTERS[18][18] ), .ZN(n1033) );
  INV_X1 U1828 ( .A(\REGISTERS[14][18] ), .ZN(n1040) );
  INV_X1 U1829 ( .A(\REGISTERS[10][18] ), .ZN(n1043) );
  INV_X1 U1830 ( .A(\REGISTERS[6][18] ), .ZN(n1046) );
  INV_X1 U1831 ( .A(\REGISTERS[2][18] ), .ZN(n1049) );
  INV_X1 U1832 ( .A(\REGISTERS[30][19] ), .ZN(n990) );
  INV_X1 U1833 ( .A(\REGISTERS[26][19] ), .ZN(n993) );
  INV_X1 U1834 ( .A(\REGISTERS[22][19] ), .ZN(n996) );
  INV_X1 U1835 ( .A(\REGISTERS[18][19] ), .ZN(n999) );
  INV_X1 U1836 ( .A(\REGISTERS[14][19] ), .ZN(n1006) );
  INV_X1 U1837 ( .A(\REGISTERS[10][19] ), .ZN(n1009) );
  INV_X1 U1838 ( .A(\REGISTERS[6][19] ), .ZN(n1012) );
  INV_X1 U1839 ( .A(\REGISTERS[2][19] ), .ZN(n1015) );
  INV_X1 U1840 ( .A(\REGISTERS[30][20] ), .ZN(n956) );
  INV_X1 U1841 ( .A(\REGISTERS[26][20] ), .ZN(n959) );
  INV_X1 U1842 ( .A(\REGISTERS[22][20] ), .ZN(n962) );
  INV_X1 U1843 ( .A(\REGISTERS[18][20] ), .ZN(n965) );
  INV_X1 U1844 ( .A(\REGISTERS[14][20] ), .ZN(n972) );
  INV_X1 U1845 ( .A(\REGISTERS[10][20] ), .ZN(n975) );
  INV_X1 U1846 ( .A(\REGISTERS[6][20] ), .ZN(n978) );
  INV_X1 U1847 ( .A(\REGISTERS[2][20] ), .ZN(n981) );
  INV_X1 U1848 ( .A(\REGISTERS[30][21] ), .ZN(n922) );
  INV_X1 U1849 ( .A(\REGISTERS[26][21] ), .ZN(n925) );
  INV_X1 U1850 ( .A(\REGISTERS[22][21] ), .ZN(n928) );
  INV_X1 U1851 ( .A(\REGISTERS[18][21] ), .ZN(n931) );
  INV_X1 U1852 ( .A(\REGISTERS[14][21] ), .ZN(n938) );
  INV_X1 U1853 ( .A(\REGISTERS[10][21] ), .ZN(n941) );
  INV_X1 U1854 ( .A(\REGISTERS[6][21] ), .ZN(n944) );
  INV_X1 U1855 ( .A(\REGISTERS[2][21] ), .ZN(n947) );
  INV_X1 U1856 ( .A(\REGISTERS[30][22] ), .ZN(n888) );
  INV_X1 U1857 ( .A(\REGISTERS[26][22] ), .ZN(n891) );
  INV_X1 U1858 ( .A(\REGISTERS[22][22] ), .ZN(n894) );
  INV_X1 U1859 ( .A(\REGISTERS[18][22] ), .ZN(n897) );
  INV_X1 U1860 ( .A(\REGISTERS[14][22] ), .ZN(n904) );
  INV_X1 U1861 ( .A(\REGISTERS[10][22] ), .ZN(n907) );
  INV_X1 U1862 ( .A(\REGISTERS[6][22] ), .ZN(n910) );
  INV_X1 U1863 ( .A(\REGISTERS[2][22] ), .ZN(n913) );
  INV_X1 U1864 ( .A(\REGISTERS[30][23] ), .ZN(n854) );
  INV_X1 U1865 ( .A(\REGISTERS[26][23] ), .ZN(n857) );
  INV_X1 U1866 ( .A(\REGISTERS[22][23] ), .ZN(n860) );
  INV_X1 U1867 ( .A(\REGISTERS[18][23] ), .ZN(n863) );
  INV_X1 U1868 ( .A(\REGISTERS[14][23] ), .ZN(n870) );
  INV_X1 U1869 ( .A(\REGISTERS[10][23] ), .ZN(n873) );
  INV_X1 U1870 ( .A(\REGISTERS[6][23] ), .ZN(n876) );
  INV_X1 U1871 ( .A(\REGISTERS[2][23] ), .ZN(n879) );
  INV_X1 U1872 ( .A(\REGISTERS[30][24] ), .ZN(n820) );
  INV_X1 U1873 ( .A(\REGISTERS[26][24] ), .ZN(n823) );
  INV_X1 U1874 ( .A(\REGISTERS[22][24] ), .ZN(n826) );
  INV_X1 U1875 ( .A(\REGISTERS[18][24] ), .ZN(n829) );
  INV_X1 U1876 ( .A(\REGISTERS[14][24] ), .ZN(n836) );
  INV_X1 U1877 ( .A(\REGISTERS[10][24] ), .ZN(n839) );
  INV_X1 U1878 ( .A(\REGISTERS[6][24] ), .ZN(n842) );
  INV_X1 U1879 ( .A(\REGISTERS[2][24] ), .ZN(n845) );
  INV_X1 U1880 ( .A(\REGISTERS[30][25] ), .ZN(n786) );
  INV_X1 U1881 ( .A(\REGISTERS[26][25] ), .ZN(n789) );
  INV_X1 U1882 ( .A(\REGISTERS[22][25] ), .ZN(n792) );
  INV_X1 U1883 ( .A(\REGISTERS[18][25] ), .ZN(n795) );
  INV_X1 U1884 ( .A(\REGISTERS[14][25] ), .ZN(n802) );
  INV_X1 U1885 ( .A(\REGISTERS[10][25] ), .ZN(n805) );
  INV_X1 U1886 ( .A(\REGISTERS[6][25] ), .ZN(n808) );
  INV_X1 U1887 ( .A(\REGISTERS[2][25] ), .ZN(n811) );
  INV_X1 U1888 ( .A(\REGISTERS[30][26] ), .ZN(n752) );
  INV_X1 U1889 ( .A(\REGISTERS[26][26] ), .ZN(n755) );
  INV_X1 U1890 ( .A(\REGISTERS[22][26] ), .ZN(n758) );
  INV_X1 U1891 ( .A(\REGISTERS[18][26] ), .ZN(n761) );
  INV_X1 U1892 ( .A(\REGISTERS[14][26] ), .ZN(n768) );
  INV_X1 U1893 ( .A(\REGISTERS[10][26] ), .ZN(n771) );
  INV_X1 U1895 ( .A(\REGISTERS[6][26] ), .ZN(n774) );
  INV_X1 U1896 ( .A(\REGISTERS[2][26] ), .ZN(n777) );
  INV_X1 U1897 ( .A(\REGISTERS[30][27] ), .ZN(n718) );
  INV_X1 U1898 ( .A(\REGISTERS[26][27] ), .ZN(n721) );
  INV_X1 U1911 ( .A(\REGISTERS[22][27] ), .ZN(n724) );
  INV_X1 U1912 ( .A(\REGISTERS[18][27] ), .ZN(n727) );
  INV_X1 U1913 ( .A(\REGISTERS[14][27] ), .ZN(n734) );
  INV_X1 U1914 ( .A(\REGISTERS[10][27] ), .ZN(n737) );
  INV_X1 U1915 ( .A(\REGISTERS[6][27] ), .ZN(n740) );
  INV_X1 U1916 ( .A(\REGISTERS[2][27] ), .ZN(n743) );
  INV_X1 U1917 ( .A(\REGISTERS[30][28] ), .ZN(n684) );
  INV_X1 U1918 ( .A(\REGISTERS[26][28] ), .ZN(n687) );
  INV_X1 U1919 ( .A(\REGISTERS[22][28] ), .ZN(n690) );
  INV_X1 U1920 ( .A(\REGISTERS[18][28] ), .ZN(n693) );
  INV_X1 U1921 ( .A(\REGISTERS[14][28] ), .ZN(n700) );
  INV_X1 U1922 ( .A(\REGISTERS[10][28] ), .ZN(n703) );
  INV_X1 U1923 ( .A(\REGISTERS[6][28] ), .ZN(n706) );
  INV_X1 U1924 ( .A(\REGISTERS[2][28] ), .ZN(n709) );
  INV_X1 U1925 ( .A(\REGISTERS[30][29] ), .ZN(n650) );
  INV_X1 U1926 ( .A(\REGISTERS[26][29] ), .ZN(n653) );
  INV_X1 U1927 ( .A(\REGISTERS[22][29] ), .ZN(n656) );
  INV_X1 U1928 ( .A(\REGISTERS[18][29] ), .ZN(n659) );
  INV_X1 U1929 ( .A(\REGISTERS[14][29] ), .ZN(n666) );
  INV_X1 U1930 ( .A(\REGISTERS[10][29] ), .ZN(n669) );
  INV_X1 U1931 ( .A(\REGISTERS[6][29] ), .ZN(n672) );
  INV_X1 U1932 ( .A(\REGISTERS[2][29] ), .ZN(n675) );
  INV_X1 U1933 ( .A(\REGISTERS[30][30] ), .ZN(n616) );
  INV_X1 U1934 ( .A(\REGISTERS[26][30] ), .ZN(n619) );
  INV_X1 U1935 ( .A(\REGISTERS[22][30] ), .ZN(n622) );
  INV_X1 U1936 ( .A(\REGISTERS[18][30] ), .ZN(n625) );
  INV_X1 U1937 ( .A(\REGISTERS[14][30] ), .ZN(n632) );
  INV_X1 U1938 ( .A(\REGISTERS[10][30] ), .ZN(n635) );
  INV_X1 U1939 ( .A(\REGISTERS[6][30] ), .ZN(n638) );
  INV_X1 U1940 ( .A(\REGISTERS[2][30] ), .ZN(n641) );
  INV_X1 U1941 ( .A(\REGISTERS[30][31] ), .ZN(n551) );
  INV_X1 U1942 ( .A(\REGISTERS[26][31] ), .ZN(n558) );
  INV_X1 U1943 ( .A(\REGISTERS[22][31] ), .ZN(n565) );
  INV_X1 U1944 ( .A(\REGISTERS[18][31] ), .ZN(n572) );
  INV_X1 U1945 ( .A(\REGISTERS[14][31] ), .ZN(n583) );
  INV_X1 U1946 ( .A(\REGISTERS[10][31] ), .ZN(n590) );
  INV_X1 U1947 ( .A(\REGISTERS[6][31] ), .ZN(n597) );
  INV_X1 U1948 ( .A(\REGISTERS[2][31] ), .ZN(n604) );
  INV_X1 U1949 ( .A(\REGISTERS[31][0] ), .ZN(n1637) );
  INV_X1 U1950 ( .A(\REGISTERS[27][0] ), .ZN(n1644) );
  INV_X1 U1951 ( .A(\REGISTERS[23][0] ), .ZN(n1650) );
  INV_X1 U1952 ( .A(\REGISTERS[19][0] ), .ZN(n1655) );
  INV_X1 U1953 ( .A(\REGISTERS[15][0] ), .ZN(n1663) );
  INV_X1 U1954 ( .A(\REGISTERS[11][0] ), .ZN(n1668) );
  INV_X1 U1955 ( .A(\REGISTERS[7][0] ), .ZN(n1671) );
  INV_X1 U1956 ( .A(\REGISTERS[3][0] ), .ZN(n1678) );
  INV_X1 U1957 ( .A(\REGISTERS[31][1] ), .ZN(n1603) );
  INV_X1 U1958 ( .A(\REGISTERS[27][1] ), .ZN(n1606) );
  INV_X1 U1959 ( .A(\REGISTERS[23][1] ), .ZN(n1609) );
  INV_X1 U1960 ( .A(\REGISTERS[19][1] ), .ZN(n1612) );
  INV_X1 U1961 ( .A(\REGISTERS[15][1] ), .ZN(n1619) );
  INV_X1 U1962 ( .A(\REGISTERS[11][1] ), .ZN(n1622) );
  INV_X1 U1963 ( .A(\REGISTERS[7][1] ), .ZN(n1625) );
  INV_X1 U1964 ( .A(\REGISTERS[3][1] ), .ZN(n1628) );
  INV_X1 U1965 ( .A(\REGISTERS[31][2] ), .ZN(n1569) );
  INV_X1 U1966 ( .A(\REGISTERS[27][2] ), .ZN(n1572) );
  INV_X1 U1967 ( .A(\REGISTERS[23][2] ), .ZN(n1575) );
  INV_X1 U1968 ( .A(\REGISTERS[19][2] ), .ZN(n1578) );
  INV_X1 U1969 ( .A(\REGISTERS[15][2] ), .ZN(n1585) );
  INV_X1 U1970 ( .A(\REGISTERS[11][2] ), .ZN(n1588) );
  INV_X1 U1971 ( .A(\REGISTERS[7][2] ), .ZN(n1591) );
  INV_X1 U1972 ( .A(\REGISTERS[3][2] ), .ZN(n1594) );
  INV_X1 U1973 ( .A(\REGISTERS[31][3] ), .ZN(n1535) );
  INV_X1 U1974 ( .A(\REGISTERS[27][3] ), .ZN(n1538) );
  INV_X1 U1975 ( .A(\REGISTERS[23][3] ), .ZN(n1541) );
  INV_X1 U1976 ( .A(\REGISTERS[19][3] ), .ZN(n1544) );
  INV_X1 U1977 ( .A(\REGISTERS[15][3] ), .ZN(n1551) );
  INV_X1 U1978 ( .A(\REGISTERS[11][3] ), .ZN(n1554) );
  INV_X1 U1979 ( .A(\REGISTERS[7][3] ), .ZN(n1557) );
  INV_X1 U1980 ( .A(\REGISTERS[3][3] ), .ZN(n1560) );
  INV_X1 U1981 ( .A(\REGISTERS[31][4] ), .ZN(n1501) );
  INV_X1 U1982 ( .A(\REGISTERS[27][4] ), .ZN(n1504) );
  INV_X1 U1983 ( .A(\REGISTERS[23][4] ), .ZN(n1507) );
  INV_X1 U1984 ( .A(\REGISTERS[19][4] ), .ZN(n1510) );
  INV_X1 U1985 ( .A(\REGISTERS[15][4] ), .ZN(n1517) );
  INV_X1 U1986 ( .A(\REGISTERS[11][4] ), .ZN(n1520) );
  INV_X1 U1987 ( .A(\REGISTERS[7][4] ), .ZN(n1523) );
  INV_X1 U1988 ( .A(\REGISTERS[3][4] ), .ZN(n1526) );
  INV_X1 U1989 ( .A(\REGISTERS[31][5] ), .ZN(n1467) );
  INV_X1 U1990 ( .A(\REGISTERS[27][5] ), .ZN(n1470) );
  INV_X1 U1991 ( .A(\REGISTERS[23][5] ), .ZN(n1473) );
  INV_X1 U1992 ( .A(\REGISTERS[19][5] ), .ZN(n1476) );
  INV_X1 U1993 ( .A(\REGISTERS[15][5] ), .ZN(n1483) );
  INV_X1 U1994 ( .A(\REGISTERS[11][5] ), .ZN(n1486) );
  INV_X1 U1995 ( .A(\REGISTERS[7][5] ), .ZN(n1489) );
  INV_X1 U1996 ( .A(\REGISTERS[3][5] ), .ZN(n1492) );
  INV_X1 U1997 ( .A(\REGISTERS[31][6] ), .ZN(n1433) );
  INV_X1 U1998 ( .A(\REGISTERS[27][6] ), .ZN(n1436) );
  INV_X1 U1999 ( .A(\REGISTERS[23][6] ), .ZN(n1439) );
  INV_X1 U2000 ( .A(\REGISTERS[19][6] ), .ZN(n1442) );
  INV_X1 U2001 ( .A(\REGISTERS[15][6] ), .ZN(n1449) );
  INV_X1 U2002 ( .A(\REGISTERS[11][6] ), .ZN(n1452) );
  INV_X1 U2003 ( .A(\REGISTERS[7][6] ), .ZN(n1455) );
  INV_X1 U2004 ( .A(\REGISTERS[3][6] ), .ZN(n1458) );
  INV_X1 U2005 ( .A(\REGISTERS[31][7] ), .ZN(n1399) );
  INV_X1 U2006 ( .A(\REGISTERS[27][7] ), .ZN(n1402) );
  INV_X1 U2007 ( .A(\REGISTERS[23][7] ), .ZN(n1405) );
  INV_X1 U2008 ( .A(\REGISTERS[19][7] ), .ZN(n1408) );
  INV_X1 U2009 ( .A(\REGISTERS[15][7] ), .ZN(n1415) );
  INV_X1 U2010 ( .A(\REGISTERS[11][7] ), .ZN(n1418) );
  INV_X1 U2011 ( .A(\REGISTERS[7][7] ), .ZN(n1421) );
  INV_X1 U2012 ( .A(\REGISTERS[3][7] ), .ZN(n1424) );
  INV_X1 U2013 ( .A(\REGISTERS[31][8] ), .ZN(n1365) );
  INV_X1 U2014 ( .A(\REGISTERS[27][8] ), .ZN(n1368) );
  INV_X1 U2015 ( .A(\REGISTERS[23][8] ), .ZN(n1371) );
  INV_X1 U2016 ( .A(\REGISTERS[19][8] ), .ZN(n1374) );
  INV_X1 U2017 ( .A(\REGISTERS[15][8] ), .ZN(n1381) );
  INV_X1 U2018 ( .A(\REGISTERS[11][8] ), .ZN(n1384) );
  INV_X1 U2019 ( .A(\REGISTERS[7][8] ), .ZN(n1387) );
  INV_X1 U2020 ( .A(\REGISTERS[3][8] ), .ZN(n1390) );
  INV_X1 U2021 ( .A(\REGISTERS[31][9] ), .ZN(n1331) );
  INV_X1 U2022 ( .A(\REGISTERS[27][9] ), .ZN(n1334) );
  INV_X1 U2023 ( .A(\REGISTERS[23][9] ), .ZN(n1337) );
  INV_X1 U2024 ( .A(\REGISTERS[19][9] ), .ZN(n1340) );
  INV_X1 U2025 ( .A(\REGISTERS[15][9] ), .ZN(n1347) );
  INV_X1 U2026 ( .A(\REGISTERS[11][9] ), .ZN(n1350) );
  INV_X1 U2027 ( .A(\REGISTERS[7][9] ), .ZN(n1353) );
  INV_X1 U2028 ( .A(\REGISTERS[3][9] ), .ZN(n1356) );
  INV_X1 U2029 ( .A(\REGISTERS[31][10] ), .ZN(n1297) );
  INV_X1 U2030 ( .A(\REGISTERS[27][10] ), .ZN(n1300) );
  INV_X1 U2031 ( .A(\REGISTERS[23][10] ), .ZN(n1303) );
  INV_X1 U2032 ( .A(\REGISTERS[19][10] ), .ZN(n1306) );
  INV_X1 U2033 ( .A(\REGISTERS[15][10] ), .ZN(n1313) );
  INV_X1 U2034 ( .A(\REGISTERS[11][10] ), .ZN(n1316) );
  INV_X1 U2035 ( .A(\REGISTERS[7][10] ), .ZN(n1319) );
  INV_X1 U2036 ( .A(\REGISTERS[3][10] ), .ZN(n1322) );
  INV_X1 U2037 ( .A(\REGISTERS[31][11] ), .ZN(n1263) );
  INV_X1 U2038 ( .A(\REGISTERS[27][11] ), .ZN(n1266) );
  INV_X1 U2039 ( .A(\REGISTERS[23][11] ), .ZN(n1269) );
  INV_X1 U2040 ( .A(\REGISTERS[19][11] ), .ZN(n1272) );
  INV_X1 U2041 ( .A(\REGISTERS[15][11] ), .ZN(n1279) );
  INV_X1 U2042 ( .A(\REGISTERS[11][11] ), .ZN(n1282) );
  INV_X1 U2043 ( .A(\REGISTERS[7][11] ), .ZN(n1285) );
  INV_X1 U2044 ( .A(\REGISTERS[3][11] ), .ZN(n1288) );
  INV_X1 U2045 ( .A(\REGISTERS[31][12] ), .ZN(n1229) );
  INV_X1 U2046 ( .A(\REGISTERS[27][12] ), .ZN(n1232) );
  INV_X1 U2047 ( .A(\REGISTERS[23][12] ), .ZN(n1235) );
  INV_X1 U2048 ( .A(\REGISTERS[19][12] ), .ZN(n1238) );
  INV_X1 U2049 ( .A(\REGISTERS[15][12] ), .ZN(n1245) );
  INV_X1 U2050 ( .A(\REGISTERS[11][12] ), .ZN(n1248) );
  INV_X1 U2051 ( .A(\REGISTERS[7][12] ), .ZN(n1251) );
  INV_X1 U2052 ( .A(\REGISTERS[3][12] ), .ZN(n1254) );
  INV_X1 U2053 ( .A(\REGISTERS[31][13] ), .ZN(n1195) );
  INV_X1 U2054 ( .A(\REGISTERS[27][13] ), .ZN(n1198) );
  INV_X1 U2055 ( .A(\REGISTERS[23][13] ), .ZN(n1201) );
  INV_X1 U2056 ( .A(\REGISTERS[19][13] ), .ZN(n1204) );
  INV_X1 U2057 ( .A(\REGISTERS[15][13] ), .ZN(n1211) );
  INV_X1 U2058 ( .A(\REGISTERS[11][13] ), .ZN(n1214) );
  INV_X1 U2059 ( .A(\REGISTERS[7][13] ), .ZN(n1217) );
  INV_X1 U2060 ( .A(\REGISTERS[3][13] ), .ZN(n1220) );
  INV_X1 U2061 ( .A(\REGISTERS[31][14] ), .ZN(n1161) );
  INV_X1 U2062 ( .A(\REGISTERS[27][14] ), .ZN(n1164) );
  INV_X1 U2063 ( .A(\REGISTERS[23][14] ), .ZN(n1167) );
  INV_X1 U2064 ( .A(\REGISTERS[19][14] ), .ZN(n1170) );
  INV_X1 U2065 ( .A(\REGISTERS[15][14] ), .ZN(n1177) );
  INV_X1 U2066 ( .A(\REGISTERS[11][14] ), .ZN(n1180) );
  INV_X1 U2067 ( .A(\REGISTERS[7][14] ), .ZN(n1183) );
  INV_X1 U2068 ( .A(\REGISTERS[3][14] ), .ZN(n1186) );
  INV_X1 U2069 ( .A(\REGISTERS[31][15] ), .ZN(n1127) );
  INV_X1 U2070 ( .A(\REGISTERS[27][15] ), .ZN(n1130) );
  INV_X1 U2071 ( .A(\REGISTERS[23][15] ), .ZN(n1133) );
  INV_X1 U2072 ( .A(\REGISTERS[19][15] ), .ZN(n1136) );
  INV_X1 U2073 ( .A(\REGISTERS[15][15] ), .ZN(n1143) );
  INV_X1 U2074 ( .A(\REGISTERS[11][15] ), .ZN(n1146) );
  INV_X1 U2075 ( .A(\REGISTERS[7][15] ), .ZN(n1149) );
  INV_X1 U2076 ( .A(\REGISTERS[3][15] ), .ZN(n1152) );
  INV_X1 U2077 ( .A(\REGISTERS[31][16] ), .ZN(n1093) );
  INV_X1 U2078 ( .A(\REGISTERS[27][16] ), .ZN(n1096) );
  INV_X1 U2079 ( .A(\REGISTERS[23][16] ), .ZN(n1099) );
  INV_X1 U2080 ( .A(\REGISTERS[19][16] ), .ZN(n1102) );
  INV_X1 U2081 ( .A(\REGISTERS[15][16] ), .ZN(n1109) );
  INV_X1 U2082 ( .A(\REGISTERS[11][16] ), .ZN(n1112) );
  INV_X1 U2083 ( .A(\REGISTERS[7][16] ), .ZN(n1115) );
  INV_X1 U2084 ( .A(\REGISTERS[3][16] ), .ZN(n1118) );
  INV_X1 U2085 ( .A(\REGISTERS[31][17] ), .ZN(n1059) );
  INV_X1 U2086 ( .A(\REGISTERS[27][17] ), .ZN(n1062) );
  INV_X1 U2087 ( .A(\REGISTERS[23][17] ), .ZN(n1065) );
  INV_X1 U2088 ( .A(\REGISTERS[19][17] ), .ZN(n1068) );
  INV_X1 U2089 ( .A(\REGISTERS[15][17] ), .ZN(n1075) );
  INV_X1 U2090 ( .A(\REGISTERS[11][17] ), .ZN(n1078) );
  INV_X1 U2091 ( .A(\REGISTERS[7][17] ), .ZN(n1081) );
  INV_X1 U2092 ( .A(\REGISTERS[3][17] ), .ZN(n1084) );
  INV_X1 U2093 ( .A(\REGISTERS[31][18] ), .ZN(n1025) );
  INV_X1 U2094 ( .A(\REGISTERS[27][18] ), .ZN(n1028) );
  INV_X1 U2095 ( .A(\REGISTERS[23][18] ), .ZN(n1031) );
  INV_X1 U2096 ( .A(\REGISTERS[19][18] ), .ZN(n1034) );
  INV_X1 U2097 ( .A(\REGISTERS[15][18] ), .ZN(n1041) );
  INV_X1 U2098 ( .A(\REGISTERS[11][18] ), .ZN(n1044) );
  INV_X1 U2099 ( .A(\REGISTERS[7][18] ), .ZN(n1047) );
  INV_X1 U2100 ( .A(\REGISTERS[3][18] ), .ZN(n1050) );
  INV_X1 U2101 ( .A(\REGISTERS[31][19] ), .ZN(n991) );
  INV_X1 U2102 ( .A(\REGISTERS[27][19] ), .ZN(n994) );
  INV_X1 U2103 ( .A(\REGISTERS[23][19] ), .ZN(n997) );
  INV_X1 U2104 ( .A(\REGISTERS[19][19] ), .ZN(n1000) );
  INV_X1 U2105 ( .A(\REGISTERS[15][19] ), .ZN(n1007) );
  INV_X1 U2106 ( .A(\REGISTERS[11][19] ), .ZN(n1010) );
  INV_X1 U2107 ( .A(\REGISTERS[7][19] ), .ZN(n1013) );
  INV_X1 U2108 ( .A(\REGISTERS[3][19] ), .ZN(n1016) );
  INV_X1 U2109 ( .A(\REGISTERS[31][20] ), .ZN(n957) );
  INV_X1 U2110 ( .A(\REGISTERS[27][20] ), .ZN(n960) );
  INV_X1 U2111 ( .A(\REGISTERS[23][20] ), .ZN(n963) );
  INV_X1 U2112 ( .A(\REGISTERS[19][20] ), .ZN(n966) );
  INV_X1 U2113 ( .A(\REGISTERS[15][20] ), .ZN(n973) );
  INV_X1 U2114 ( .A(\REGISTERS[11][20] ), .ZN(n976) );
  INV_X1 U2115 ( .A(\REGISTERS[7][20] ), .ZN(n979) );
  INV_X1 U2116 ( .A(\REGISTERS[3][20] ), .ZN(n982) );
  INV_X1 U2117 ( .A(\REGISTERS[31][21] ), .ZN(n923) );
  INV_X1 U2118 ( .A(\REGISTERS[27][21] ), .ZN(n926) );
  INV_X1 U2119 ( .A(\REGISTERS[23][21] ), .ZN(n929) );
  INV_X1 U2120 ( .A(\REGISTERS[19][21] ), .ZN(n932) );
  INV_X1 U2121 ( .A(\REGISTERS[15][21] ), .ZN(n939) );
  INV_X1 U2122 ( .A(\REGISTERS[11][21] ), .ZN(n942) );
  INV_X1 U2123 ( .A(\REGISTERS[7][21] ), .ZN(n945) );
  INV_X1 U2124 ( .A(\REGISTERS[3][21] ), .ZN(n948) );
  INV_X1 U2125 ( .A(\REGISTERS[31][22] ), .ZN(n889) );
  INV_X1 U2126 ( .A(\REGISTERS[27][22] ), .ZN(n892) );
  INV_X1 U2127 ( .A(\REGISTERS[23][22] ), .ZN(n895) );
  INV_X1 U2128 ( .A(\REGISTERS[19][22] ), .ZN(n898) );
  INV_X1 U2129 ( .A(\REGISTERS[15][22] ), .ZN(n905) );
  INV_X1 U2130 ( .A(\REGISTERS[11][22] ), .ZN(n908) );
  INV_X1 U2131 ( .A(\REGISTERS[7][22] ), .ZN(n911) );
  INV_X1 U2132 ( .A(\REGISTERS[3][22] ), .ZN(n914) );
  INV_X1 U2133 ( .A(\REGISTERS[31][23] ), .ZN(n855) );
  INV_X1 U2134 ( .A(\REGISTERS[27][23] ), .ZN(n858) );
  INV_X1 U2135 ( .A(\REGISTERS[23][23] ), .ZN(n861) );
  INV_X1 U2136 ( .A(\REGISTERS[19][23] ), .ZN(n864) );
  INV_X1 U2137 ( .A(\REGISTERS[15][23] ), .ZN(n871) );
  INV_X1 U2138 ( .A(\REGISTERS[11][23] ), .ZN(n874) );
  INV_X1 U2139 ( .A(\REGISTERS[7][23] ), .ZN(n877) );
  INV_X1 U2140 ( .A(\REGISTERS[3][23] ), .ZN(n880) );
  INV_X1 U2141 ( .A(\REGISTERS[31][24] ), .ZN(n821) );
  INV_X1 U2142 ( .A(\REGISTERS[27][24] ), .ZN(n824) );
  INV_X1 U2143 ( .A(\REGISTERS[23][24] ), .ZN(n827) );
  INV_X1 U2144 ( .A(\REGISTERS[19][24] ), .ZN(n830) );
  INV_X1 U2145 ( .A(\REGISTERS[15][24] ), .ZN(n837) );
  INV_X1 U2146 ( .A(\REGISTERS[11][24] ), .ZN(n840) );
  INV_X1 U2147 ( .A(\REGISTERS[7][24] ), .ZN(n843) );
  INV_X1 U2148 ( .A(\REGISTERS[3][24] ), .ZN(n846) );
  INV_X1 U2149 ( .A(\REGISTERS[31][25] ), .ZN(n787) );
  INV_X1 U2150 ( .A(\REGISTERS[27][25] ), .ZN(n790) );
  INV_X1 U2151 ( .A(\REGISTERS[23][25] ), .ZN(n793) );
  INV_X1 U2152 ( .A(\REGISTERS[19][25] ), .ZN(n796) );
  INV_X1 U2153 ( .A(\REGISTERS[15][25] ), .ZN(n803) );
  INV_X1 U2154 ( .A(\REGISTERS[11][25] ), .ZN(n806) );
  INV_X1 U2155 ( .A(\REGISTERS[7][25] ), .ZN(n809) );
  INV_X1 U2156 ( .A(\REGISTERS[3][25] ), .ZN(n812) );
  INV_X1 U2157 ( .A(\REGISTERS[31][26] ), .ZN(n753) );
  INV_X1 U2158 ( .A(\REGISTERS[27][26] ), .ZN(n756) );
  INV_X1 U2159 ( .A(\REGISTERS[23][26] ), .ZN(n759) );
  INV_X1 U2160 ( .A(\REGISTERS[19][26] ), .ZN(n762) );
  INV_X1 U2161 ( .A(\REGISTERS[15][26] ), .ZN(n769) );
  INV_X1 U2162 ( .A(\REGISTERS[11][26] ), .ZN(n772) );
  INV_X1 U2163 ( .A(\REGISTERS[7][26] ), .ZN(n775) );
  INV_X1 U2164 ( .A(\REGISTERS[3][26] ), .ZN(n778) );
  INV_X1 U2165 ( .A(\REGISTERS[31][27] ), .ZN(n719) );
  INV_X1 U2166 ( .A(\REGISTERS[27][27] ), .ZN(n722) );
  INV_X1 U2167 ( .A(\REGISTERS[23][27] ), .ZN(n725) );
  INV_X1 U2168 ( .A(\REGISTERS[19][27] ), .ZN(n728) );
  INV_X1 U2169 ( .A(\REGISTERS[15][27] ), .ZN(n735) );
  INV_X1 U2170 ( .A(\REGISTERS[11][27] ), .ZN(n738) );
  INV_X1 U2171 ( .A(\REGISTERS[7][27] ), .ZN(n741) );
  INV_X1 U2172 ( .A(\REGISTERS[3][27] ), .ZN(n744) );
  INV_X1 U2173 ( .A(\REGISTERS[31][28] ), .ZN(n685) );
  INV_X1 U2174 ( .A(\REGISTERS[27][28] ), .ZN(n688) );
  INV_X1 U2175 ( .A(\REGISTERS[23][28] ), .ZN(n691) );
  INV_X1 U2176 ( .A(\REGISTERS[19][28] ), .ZN(n694) );
  INV_X1 U2177 ( .A(\REGISTERS[15][28] ), .ZN(n701) );
  INV_X1 U2178 ( .A(\REGISTERS[11][28] ), .ZN(n704) );
  INV_X1 U2179 ( .A(\REGISTERS[7][28] ), .ZN(n707) );
  INV_X1 U2180 ( .A(\REGISTERS[3][28] ), .ZN(n710) );
  INV_X1 U2181 ( .A(\REGISTERS[31][29] ), .ZN(n651) );
  INV_X1 U2182 ( .A(\REGISTERS[27][29] ), .ZN(n654) );
  INV_X1 U2183 ( .A(\REGISTERS[23][29] ), .ZN(n657) );
  INV_X1 U2184 ( .A(\REGISTERS[19][29] ), .ZN(n660) );
  INV_X1 U2185 ( .A(\REGISTERS[15][29] ), .ZN(n667) );
  INV_X1 U2186 ( .A(\REGISTERS[11][29] ), .ZN(n670) );
  INV_X1 U2187 ( .A(\REGISTERS[7][29] ), .ZN(n673) );
  INV_X1 U2188 ( .A(\REGISTERS[3][29] ), .ZN(n676) );
  INV_X1 U2189 ( .A(\REGISTERS[31][30] ), .ZN(n617) );
  INV_X1 U2190 ( .A(\REGISTERS[27][30] ), .ZN(n620) );
  INV_X1 U2191 ( .A(\REGISTERS[23][30] ), .ZN(n623) );
  INV_X1 U2192 ( .A(\REGISTERS[19][30] ), .ZN(n626) );
  INV_X1 U2193 ( .A(\REGISTERS[15][30] ), .ZN(n633) );
  INV_X1 U2194 ( .A(\REGISTERS[11][30] ), .ZN(n636) );
  INV_X1 U2195 ( .A(\REGISTERS[7][30] ), .ZN(n639) );
  INV_X1 U2196 ( .A(\REGISTERS[3][30] ), .ZN(n642) );
  INV_X1 U2197 ( .A(\REGISTERS[31][31] ), .ZN(n553) );
  INV_X1 U2198 ( .A(\REGISTERS[27][31] ), .ZN(n560) );
  INV_X1 U2199 ( .A(\REGISTERS[23][31] ), .ZN(n567) );
  INV_X1 U2200 ( .A(\REGISTERS[19][31] ), .ZN(n574) );
  INV_X1 U2201 ( .A(\REGISTERS[15][31] ), .ZN(n585) );
  INV_X1 U2202 ( .A(\REGISTERS[11][31] ), .ZN(n592) );
  INV_X1 U2203 ( .A(\REGISTERS[7][31] ), .ZN(n599) );
  INV_X1 U2204 ( .A(\REGISTERS[3][31] ), .ZN(n606) );
  INV_X1 U2205 ( .A(ADD_RD1[1]), .ZN(n2301) );
  CLKBUF_X1 U2206 ( .A(n4612), .Z(n4812) );
  CLKBUF_X1 U2207 ( .A(n4612), .Z(n4813) );
  CLKBUF_X1 U2208 ( .A(n4612), .Z(n4814) );
  CLKBUF_X1 U2209 ( .A(n4612), .Z(n4815) );
  CLKBUF_X1 U2210 ( .A(n4608), .Z(n4816) );
  CLKBUF_X1 U2211 ( .A(n4608), .Z(n4817) );
  CLKBUF_X1 U2212 ( .A(n4608), .Z(n4818) );
  CLKBUF_X1 U2213 ( .A(n4608), .Z(n4819) );
  CLKBUF_X1 U2214 ( .A(n4604), .Z(n4820) );
  CLKBUF_X1 U2215 ( .A(n4604), .Z(n4821) );
  CLKBUF_X1 U2216 ( .A(n4604), .Z(n4822) );
  CLKBUF_X1 U2217 ( .A(n4604), .Z(n4823) );
  CLKBUF_X1 U2218 ( .A(n4600), .Z(n4824) );
  CLKBUF_X1 U2219 ( .A(n4600), .Z(n4825) );
  CLKBUF_X1 U2220 ( .A(n4600), .Z(n4826) );
  CLKBUF_X1 U2221 ( .A(n4600), .Z(n4827) );
  CLKBUF_X1 U2222 ( .A(n4596), .Z(n4828) );
  CLKBUF_X1 U2223 ( .A(n4596), .Z(n4829) );
  CLKBUF_X1 U2224 ( .A(n4596), .Z(n4830) );
  CLKBUF_X1 U2225 ( .A(n4596), .Z(n4831) );
  CLKBUF_X1 U2226 ( .A(n4592), .Z(n4832) );
  CLKBUF_X1 U2227 ( .A(n4592), .Z(n4833) );
  CLKBUF_X1 U2228 ( .A(n4592), .Z(n4834) );
  CLKBUF_X1 U2229 ( .A(n4592), .Z(n4835) );
  CLKBUF_X1 U2230 ( .A(n4588), .Z(n4836) );
  CLKBUF_X1 U2231 ( .A(n4588), .Z(n4837) );
  CLKBUF_X1 U2232 ( .A(n4588), .Z(n4838) );
  CLKBUF_X1 U2233 ( .A(n4588), .Z(n4839) );
  CLKBUF_X1 U2234 ( .A(n4584), .Z(n4840) );
  CLKBUF_X1 U2235 ( .A(n4584), .Z(n4841) );
  CLKBUF_X1 U2236 ( .A(n4584), .Z(n4842) );
  CLKBUF_X1 U2237 ( .A(n4584), .Z(n4843) );
  CLKBUF_X1 U2238 ( .A(n4580), .Z(n4844) );
  CLKBUF_X1 U2239 ( .A(n4580), .Z(n4845) );
  CLKBUF_X1 U2240 ( .A(n4580), .Z(n4846) );
  CLKBUF_X1 U2241 ( .A(n4580), .Z(n4847) );
  CLKBUF_X1 U2242 ( .A(n4576), .Z(n4848) );
  CLKBUF_X1 U2243 ( .A(n4576), .Z(n4849) );
  CLKBUF_X1 U2244 ( .A(n4576), .Z(n4850) );
  CLKBUF_X1 U2245 ( .A(n4576), .Z(n4851) );
  CLKBUF_X1 U2246 ( .A(n4572), .Z(n4852) );
  CLKBUF_X1 U2247 ( .A(n4572), .Z(n4853) );
  CLKBUF_X1 U2248 ( .A(n4572), .Z(n4854) );
  CLKBUF_X1 U2249 ( .A(n4572), .Z(n4855) );
  CLKBUF_X1 U2250 ( .A(n4568), .Z(n4856) );
  CLKBUF_X1 U2251 ( .A(n4568), .Z(n4857) );
  CLKBUF_X1 U2252 ( .A(n4568), .Z(n4858) );
  CLKBUF_X1 U2253 ( .A(n4568), .Z(n4859) );
  CLKBUF_X1 U2254 ( .A(n4564), .Z(n4860) );
  CLKBUF_X1 U2255 ( .A(n4564), .Z(n4861) );
  CLKBUF_X1 U2256 ( .A(n4564), .Z(n4862) );
  CLKBUF_X1 U2257 ( .A(n4564), .Z(n4863) );
  CLKBUF_X1 U2258 ( .A(n4560), .Z(n4864) );
  CLKBUF_X1 U2259 ( .A(n4560), .Z(n4865) );
  CLKBUF_X1 U2260 ( .A(n4560), .Z(n4866) );
  CLKBUF_X1 U2261 ( .A(n4560), .Z(n4867) );
  CLKBUF_X1 U2262 ( .A(n4556), .Z(n4868) );
  CLKBUF_X1 U2263 ( .A(n4556), .Z(n4869) );
  CLKBUF_X1 U2264 ( .A(n4556), .Z(n4870) );
  CLKBUF_X1 U2265 ( .A(n4556), .Z(n4871) );
  CLKBUF_X1 U2266 ( .A(n4552), .Z(n4872) );
  CLKBUF_X1 U2267 ( .A(n4552), .Z(n4873) );
  CLKBUF_X1 U2268 ( .A(n4552), .Z(n4874) );
  CLKBUF_X1 U2269 ( .A(n4552), .Z(n4875) );
  CLKBUF_X1 U2270 ( .A(n4548), .Z(n4876) );
  CLKBUF_X1 U2271 ( .A(n4548), .Z(n4877) );
  CLKBUF_X1 U2272 ( .A(n4548), .Z(n4878) );
  CLKBUF_X1 U2273 ( .A(n4548), .Z(n4879) );
  CLKBUF_X1 U2274 ( .A(n4544), .Z(n4880) );
  CLKBUF_X1 U2275 ( .A(n4544), .Z(n4881) );
  CLKBUF_X1 U2276 ( .A(n4544), .Z(n4882) );
  CLKBUF_X1 U2277 ( .A(n4544), .Z(n4883) );
  CLKBUF_X1 U2278 ( .A(n4540), .Z(n4884) );
  CLKBUF_X1 U2279 ( .A(n4540), .Z(n4885) );
  CLKBUF_X1 U2280 ( .A(n4540), .Z(n4886) );
  CLKBUF_X1 U2281 ( .A(n4540), .Z(n4887) );
  CLKBUF_X1 U2282 ( .A(n4536), .Z(n4888) );
  CLKBUF_X1 U2283 ( .A(n4536), .Z(n4889) );
  CLKBUF_X1 U2284 ( .A(n4536), .Z(n4890) );
  CLKBUF_X1 U2285 ( .A(n4536), .Z(n4891) );
  CLKBUF_X1 U2286 ( .A(n4532), .Z(n4892) );
  CLKBUF_X1 U2287 ( .A(n4532), .Z(n4893) );
  CLKBUF_X1 U2288 ( .A(n4532), .Z(n4894) );
  CLKBUF_X1 U2289 ( .A(n4532), .Z(n4895) );
  CLKBUF_X1 U2290 ( .A(n4528), .Z(n4896) );
  CLKBUF_X1 U2291 ( .A(n4528), .Z(n4897) );
  CLKBUF_X1 U2292 ( .A(n4528), .Z(n4898) );
  CLKBUF_X1 U2293 ( .A(n4528), .Z(n4899) );
  CLKBUF_X1 U2294 ( .A(n4524), .Z(n4900) );
  CLKBUF_X1 U2295 ( .A(n4524), .Z(n4901) );
  CLKBUF_X1 U2296 ( .A(n4524), .Z(n4902) );
  CLKBUF_X1 U2297 ( .A(n4524), .Z(n4903) );
  CLKBUF_X1 U2298 ( .A(n4520), .Z(n4904) );
  CLKBUF_X1 U2299 ( .A(n4520), .Z(n4905) );
  CLKBUF_X1 U2300 ( .A(n4520), .Z(n4906) );
  CLKBUF_X1 U2301 ( .A(n4520), .Z(n4907) );
  CLKBUF_X1 U2302 ( .A(n4516), .Z(n4908) );
  CLKBUF_X1 U2303 ( .A(n4516), .Z(n4909) );
  CLKBUF_X1 U2304 ( .A(n4516), .Z(n4910) );
  CLKBUF_X1 U2305 ( .A(n4516), .Z(n4911) );
  CLKBUF_X1 U2306 ( .A(n4512), .Z(n4912) );
  CLKBUF_X1 U2307 ( .A(n4512), .Z(n4913) );
  CLKBUF_X1 U2308 ( .A(n4512), .Z(n4914) );
  CLKBUF_X1 U2309 ( .A(n4512), .Z(n4915) );
  CLKBUF_X1 U2310 ( .A(n4508), .Z(n4916) );
  CLKBUF_X1 U2311 ( .A(n4508), .Z(n4917) );
  CLKBUF_X1 U2312 ( .A(n4508), .Z(n4918) );
  CLKBUF_X1 U2313 ( .A(n4508), .Z(n4919) );
  CLKBUF_X1 U2314 ( .A(n4504), .Z(n4920) );
  CLKBUF_X1 U2315 ( .A(n4504), .Z(n4921) );
  CLKBUF_X1 U2316 ( .A(n4504), .Z(n4922) );
  CLKBUF_X1 U2317 ( .A(n4504), .Z(n4923) );
  CLKBUF_X1 U2318 ( .A(n4500), .Z(n4924) );
  CLKBUF_X1 U2319 ( .A(n4500), .Z(n4925) );
  CLKBUF_X1 U2320 ( .A(n4500), .Z(n4926) );
  CLKBUF_X1 U2321 ( .A(n4500), .Z(n4927) );
  CLKBUF_X1 U2322 ( .A(n4496), .Z(n4928) );
  CLKBUF_X1 U2323 ( .A(n4496), .Z(n4929) );
  CLKBUF_X1 U2324 ( .A(n4496), .Z(n4930) );
  CLKBUF_X1 U2325 ( .A(n4496), .Z(n4931) );
  CLKBUF_X1 U2326 ( .A(n4492), .Z(n4932) );
  CLKBUF_X1 U2327 ( .A(n4492), .Z(n4933) );
  CLKBUF_X1 U2328 ( .A(n4492), .Z(n4934) );
  CLKBUF_X1 U2329 ( .A(n4492), .Z(n4935) );
  CLKBUF_X1 U2330 ( .A(n4488), .Z(n4936) );
  CLKBUF_X1 U2331 ( .A(n4488), .Z(n4937) );
  CLKBUF_X1 U2332 ( .A(n4488), .Z(n4938) );
  CLKBUF_X1 U2333 ( .A(n4488), .Z(n4939) );
  CLKBUF_X1 U2334 ( .A(n4484), .Z(n4940) );
  CLKBUF_X1 U2335 ( .A(n4484), .Z(n4941) );
  CLKBUF_X1 U2336 ( .A(n4484), .Z(n4942) );
  CLKBUF_X1 U2337 ( .A(n4484), .Z(n4943) );
  CLKBUF_X1 U2338 ( .A(n4480), .Z(n4947) );
  CLKBUF_X1 U2339 ( .A(n4476), .Z(n4951) );
  CLKBUF_X1 U2340 ( .A(n4472), .Z(n4955) );
  CLKBUF_X1 U2341 ( .A(n4468), .Z(n4959) );
  CLKBUF_X1 U2342 ( .A(n4464), .Z(n4963) );
  CLKBUF_X1 U2343 ( .A(n4460), .Z(n4967) );
  CLKBUF_X1 U2344 ( .A(n4456), .Z(n4971) );
  CLKBUF_X1 U2345 ( .A(n4452), .Z(n4975) );
  CLKBUF_X1 U2346 ( .A(n4448), .Z(n4979) );
  CLKBUF_X1 U2347 ( .A(n4444), .Z(n4983) );
  CLKBUF_X1 U2348 ( .A(n4440), .Z(n4987) );
  CLKBUF_X1 U2349 ( .A(n4436), .Z(n4991) );
  CLKBUF_X1 U2350 ( .A(n4432), .Z(n4995) );
  CLKBUF_X1 U2351 ( .A(n4428), .Z(n4999) );
  CLKBUF_X1 U2352 ( .A(n4424), .Z(n5003) );
  CLKBUF_X1 U2353 ( .A(n4420), .Z(n5007) );
  CLKBUF_X1 U2354 ( .A(n4416), .Z(n5011) );
  CLKBUF_X1 U2355 ( .A(n4412), .Z(n5015) );
  CLKBUF_X1 U2356 ( .A(n4408), .Z(n5019) );
  CLKBUF_X1 U2357 ( .A(n4404), .Z(n5023) );
  CLKBUF_X1 U2358 ( .A(n4400), .Z(n5027) );
  CLKBUF_X1 U2359 ( .A(n4396), .Z(n5031) );
  CLKBUF_X1 U2360 ( .A(n4392), .Z(n5035) );
  CLKBUF_X1 U2361 ( .A(n4388), .Z(n5039) );
  CLKBUF_X1 U2362 ( .A(n4384), .Z(n5043) );
  CLKBUF_X1 U2363 ( .A(n4380), .Z(n5047) );
  CLKBUF_X1 U2364 ( .A(n4376), .Z(n5051) );
  CLKBUF_X1 U2365 ( .A(n4372), .Z(n5055) );
  CLKBUF_X1 U2366 ( .A(n4368), .Z(n5059) );
  CLKBUF_X1 U2367 ( .A(n4364), .Z(n5063) );
  CLKBUF_X1 U2368 ( .A(n4360), .Z(n5067) );
  CLKBUF_X1 U2369 ( .A(n4356), .Z(n5068) );
  CLKBUF_X1 U2370 ( .A(n4356), .Z(n5069) );
  CLKBUF_X1 U2371 ( .A(n4356), .Z(n5070) );
  CLKBUF_X1 U2372 ( .A(n4356), .Z(n5071) );
  CLKBUF_X1 U2373 ( .A(n4352), .Z(n5075) );
endmodule


module DLX_IR_SIZE32_PC_SIZE32_DW01_add_1 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \A[1] , \A[0] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , n1;
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];
  assign \carry[3]  = A[2];

  XOR2_X1 U3 ( .A(A[30]), .B(\carry[30] ), .Z(SUM[30]) );
  XOR2_X1 U5 ( .A(A[29]), .B(\carry[29] ), .Z(SUM[29]) );
  XOR2_X1 U7 ( .A(A[28]), .B(\carry[28] ), .Z(SUM[28]) );
  XOR2_X1 U9 ( .A(A[27]), .B(\carry[27] ), .Z(SUM[27]) );
  XOR2_X1 U11 ( .A(A[26]), .B(\carry[26] ), .Z(SUM[26]) );
  XOR2_X1 U13 ( .A(A[25]), .B(\carry[25] ), .Z(SUM[25]) );
  XOR2_X1 U15 ( .A(A[24]), .B(\carry[24] ), .Z(SUM[24]) );
  XOR2_X1 U17 ( .A(A[23]), .B(\carry[23] ), .Z(SUM[23]) );
  XOR2_X1 U19 ( .A(A[22]), .B(\carry[22] ), .Z(SUM[22]) );
  XOR2_X1 U21 ( .A(A[21]), .B(\carry[21] ), .Z(SUM[21]) );
  XOR2_X1 U23 ( .A(A[20]), .B(\carry[20] ), .Z(SUM[20]) );
  XOR2_X1 U25 ( .A(A[19]), .B(\carry[19] ), .Z(SUM[19]) );
  XOR2_X1 U27 ( .A(A[18]), .B(\carry[18] ), .Z(SUM[18]) );
  XOR2_X1 U29 ( .A(A[17]), .B(\carry[17] ), .Z(SUM[17]) );
  XOR2_X1 U31 ( .A(A[16]), .B(\carry[16] ), .Z(SUM[16]) );
  XOR2_X1 U33 ( .A(A[15]), .B(\carry[15] ), .Z(SUM[15]) );
  XOR2_X1 U35 ( .A(A[14]), .B(\carry[14] ), .Z(SUM[14]) );
  XOR2_X1 U37 ( .A(A[13]), .B(\carry[13] ), .Z(SUM[13]) );
  XOR2_X1 U39 ( .A(A[12]), .B(\carry[12] ), .Z(SUM[12]) );
  XOR2_X1 U41 ( .A(A[11]), .B(\carry[11] ), .Z(SUM[11]) );
  XOR2_X1 U43 ( .A(A[10]), .B(\carry[10] ), .Z(SUM[10]) );
  XOR2_X1 U45 ( .A(A[9]), .B(\carry[9] ), .Z(SUM[9]) );
  XOR2_X1 U47 ( .A(A[8]), .B(\carry[8] ), .Z(SUM[8]) );
  XOR2_X1 U49 ( .A(A[7]), .B(\carry[7] ), .Z(SUM[7]) );
  XOR2_X1 U51 ( .A(A[6]), .B(\carry[6] ), .Z(SUM[6]) );
  XOR2_X1 U53 ( .A(A[5]), .B(\carry[5] ), .Z(SUM[5]) );
  XOR2_X1 U55 ( .A(A[4]), .B(\carry[4] ), .Z(SUM[4]) );
  XOR2_X1 U57 ( .A(A[3]), .B(\carry[3] ), .Z(SUM[3]) );
  XNOR2_X1 U1 ( .A(A[31]), .B(n1), .ZN(SUM[31]) );
  NAND2_X1 U2 ( .A1(\carry[30] ), .A2(A[30]), .ZN(n1) );
  AND2_X1 U4 ( .A1(\carry[29] ), .A2(A[29]), .ZN(\carry[30] ) );
  AND2_X1 U6 ( .A1(\carry[3] ), .A2(A[3]), .ZN(\carry[4] ) );
  AND2_X1 U8 ( .A1(\carry[4] ), .A2(A[4]), .ZN(\carry[5] ) );
  AND2_X1 U10 ( .A1(\carry[5] ), .A2(A[5]), .ZN(\carry[6] ) );
  AND2_X1 U12 ( .A1(\carry[6] ), .A2(A[6]), .ZN(\carry[7] ) );
  AND2_X1 U14 ( .A1(\carry[7] ), .A2(A[7]), .ZN(\carry[8] ) );
  AND2_X1 U16 ( .A1(\carry[8] ), .A2(A[8]), .ZN(\carry[9] ) );
  AND2_X1 U18 ( .A1(\carry[9] ), .A2(A[9]), .ZN(\carry[10] ) );
  AND2_X1 U20 ( .A1(\carry[10] ), .A2(A[10]), .ZN(\carry[11] ) );
  AND2_X1 U22 ( .A1(\carry[11] ), .A2(A[11]), .ZN(\carry[12] ) );
  AND2_X1 U24 ( .A1(\carry[12] ), .A2(A[12]), .ZN(\carry[13] ) );
  AND2_X1 U26 ( .A1(\carry[13] ), .A2(A[13]), .ZN(\carry[14] ) );
  AND2_X1 U28 ( .A1(\carry[14] ), .A2(A[14]), .ZN(\carry[15] ) );
  AND2_X1 U30 ( .A1(\carry[15] ), .A2(A[15]), .ZN(\carry[16] ) );
  AND2_X1 U32 ( .A1(\carry[16] ), .A2(A[16]), .ZN(\carry[17] ) );
  AND2_X1 U34 ( .A1(\carry[17] ), .A2(A[17]), .ZN(\carry[18] ) );
  AND2_X1 U36 ( .A1(\carry[18] ), .A2(A[18]), .ZN(\carry[19] ) );
  AND2_X1 U38 ( .A1(\carry[19] ), .A2(A[19]), .ZN(\carry[20] ) );
  AND2_X1 U40 ( .A1(\carry[20] ), .A2(A[20]), .ZN(\carry[21] ) );
  AND2_X1 U42 ( .A1(\carry[21] ), .A2(A[21]), .ZN(\carry[22] ) );
  AND2_X1 U44 ( .A1(\carry[22] ), .A2(A[22]), .ZN(\carry[23] ) );
  AND2_X1 U46 ( .A1(\carry[23] ), .A2(A[23]), .ZN(\carry[24] ) );
  AND2_X1 U48 ( .A1(\carry[24] ), .A2(A[24]), .ZN(\carry[25] ) );
  AND2_X1 U50 ( .A1(\carry[25] ), .A2(A[25]), .ZN(\carry[26] ) );
  AND2_X1 U52 ( .A1(\carry[26] ), .A2(A[26]), .ZN(\carry[27] ) );
  AND2_X1 U54 ( .A1(\carry[27] ), .A2(A[27]), .ZN(\carry[28] ) );
  AND2_X1 U56 ( .A1(\carry[28] ), .A2(A[28]), .ZN(\carry[29] ) );
  INV_X1 U58 ( .A(\carry[3] ), .ZN(SUM[2]) );
endmodule


module DLX_IR_SIZE32_PC_SIZE32_DW01_add_0 ( A, B, CI, SUM, CO );
  input [31:0] A;
  input [31:0] B;
  output [31:0] SUM;
  input CI;
  output CO;
  wire   \carry[31] , \carry[30] , \carry[29] , \carry[28] , \carry[27] ,
         \carry[26] , \carry[25] , \carry[24] , \carry[23] , \carry[22] ,
         \carry[21] , \carry[20] , \carry[19] , \carry[18] , \carry[17] ,
         \carry[16] , \carry[15] , \carry[14] , \carry[13] , \carry[12] ,
         \carry[11] , \carry[10] , \carry[9] , \carry[8] , \carry[7] ,
         \carry[6] , \carry[5] , \carry[4] , \carry[3] , \carry[2] ,
         \carry[1] ;

  FA_X1 U1_31 ( .A(A[31]), .B(B[31]), .CI(\carry[31] ), .S(SUM[31]) );
  FA_X1 U1_30 ( .A(A[30]), .B(B[30]), .CI(\carry[30] ), .CO(\carry[31] ), .S(
        SUM[30]) );
  FA_X1 U1_29 ( .A(A[29]), .B(B[29]), .CI(\carry[29] ), .CO(\carry[30] ), .S(
        SUM[29]) );
  FA_X1 U1_28 ( .A(A[28]), .B(B[28]), .CI(\carry[28] ), .CO(\carry[29] ), .S(
        SUM[28]) );
  FA_X1 U1_27 ( .A(A[27]), .B(B[27]), .CI(\carry[27] ), .CO(\carry[28] ), .S(
        SUM[27]) );
  FA_X1 U1_26 ( .A(A[26]), .B(B[26]), .CI(\carry[26] ), .CO(\carry[27] ), .S(
        SUM[26]) );
  FA_X1 U1_25 ( .A(A[25]), .B(B[25]), .CI(\carry[25] ), .CO(\carry[26] ), .S(
        SUM[25]) );
  FA_X1 U1_24 ( .A(A[24]), .B(B[24]), .CI(\carry[24] ), .CO(\carry[25] ), .S(
        SUM[24]) );
  FA_X1 U1_23 ( .A(A[23]), .B(B[23]), .CI(\carry[23] ), .CO(\carry[24] ), .S(
        SUM[23]) );
  FA_X1 U1_22 ( .A(A[22]), .B(B[22]), .CI(\carry[22] ), .CO(\carry[23] ), .S(
        SUM[22]) );
  FA_X1 U1_21 ( .A(A[21]), .B(B[21]), .CI(\carry[21] ), .CO(\carry[22] ), .S(
        SUM[21]) );
  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(\carry[20] ), .CO(\carry[21] ), .S(
        SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(\carry[19] ), .CO(\carry[20] ), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(\carry[18] ), .CO(\carry[19] ), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(\carry[17] ), .CO(\carry[18] ), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(\carry[16] ), .CO(\carry[17] ), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(\carry[15] ), .CO(\carry[16] ), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(\carry[14] ), .CO(\carry[15] ), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(\carry[13] ), .CO(\carry[14] ), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(\carry[12] ), .CO(\carry[13] ), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(\carry[11] ), .CO(\carry[12] ), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(\carry[10] ), .CO(\carry[11] ), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(\carry[9] ), .CO(\carry[10] ), .S(
        SUM[9]) );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(\carry[8] ), .CO(\carry[9] ), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(\carry[7] ), .CO(\carry[8] ), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(\carry[6] ), .CO(\carry[7] ), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(\carry[5] ), .CO(\carry[6] ), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(\carry[4] ), .CO(\carry[5] ), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(\carry[3] ), .CO(\carry[4] ), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(\carry[2] ), .CO(\carry[3] ), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(\carry[1] ), .CO(\carry[2] ), .S(SUM[1]) );
  XOR2_X1 U2 ( .A(B[0]), .B(A[0]), .Z(SUM[0]) );
  AND2_X1 U1 ( .A1(A[0]), .A2(B[0]), .ZN(\carry[1] ) );
endmodule



    module CU_HDW_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE21 ( 
        Clk, Rst, IR_IN, flush, IR_LATCH_EN, NPC1_LATCH_EN, NPC2_LATCH_EN, 
        RegA_LATCH_EN, RegB_LATCH_EN, RegAluOpCodeGen_EN, RegIMM_LATCH_EN, 
        Reg_RD1_EN, RD1, RD2, B2_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
        RETURN_REG_EN, Reg_RD2_EN, DRAM_WE, ALU_OUT2_SEL, LMD_LATCH_EN, 
        Alu_outreg2_en, JUMP_en, PC_LATCH_EN, Reg_RD3_EN, write_stop_if_branch, 
        WB_MUX_SEL, RF_WE, WB_MUX_ADD_SEL, WR );
  input [31:0] IR_IN;
  input Clk, Rst, flush;
  output IR_LATCH_EN, NPC1_LATCH_EN, NPC2_LATCH_EN, RegA_LATCH_EN,
         RegB_LATCH_EN, RegAluOpCodeGen_EN, RegIMM_LATCH_EN, Reg_RD1_EN, RD1,
         RD2, B2_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, RETURN_REG_EN,
         Reg_RD2_EN, DRAM_WE, ALU_OUT2_SEL, LMD_LATCH_EN, Alu_outreg2_en,
         JUMP_en, PC_LATCH_EN, Reg_RD3_EN, write_stop_if_branch, WB_MUX_SEL,
         RF_WE, WB_MUX_ADD_SEL, WR;
  wire   IR_IN_31, IR_IN_30, IR_IN_29, IR_IN_28, IR_IN_27, IR_IN_26,
         RegAluOpCodeGen_EN, N442, n42, n48, n54, n60, n65, n70, n75, n80, n85,
         n90, n95, n99, n103, n107, n111, n115, n118, n121, n124, n127, n129,
         n131, n133, n135, n137, n139, n141, n143, n145, n147, n149, n151,
         n153, n155, n157, n159, n161, n163, n165, n167, n169, RETURN_REG_EN,
         n209, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n40, n41, n46, n47, n52, n53, n55, n58, n59, n63,
         n64, n68, n69, n73, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221;
  wire   [20:0] cw;
  wire   [10:0] cw3;
  wire   [3:0] cw4;
  tri   Reg_RD1_EN;
  tri   [19:0] cw1;
  tri   [15:0] cw2;
  tri   NPC1_LATCH_EN;
  tri   RegIMM_LATCH_EN;
  tri   RD1;
  tri   RD2;
  assign IR_IN_31 = IR_IN[31];
  assign IR_IN_30 = IR_IN[30];
  assign IR_IN_29 = IR_IN[29];
  assign IR_IN_28 = IR_IN[28];
  assign IR_IN_27 = IR_IN[27];
  assign IR_IN_26 = IR_IN[26];
  assign NPC2_LATCH_EN = RegAluOpCodeGen_EN;
  assign B2_LATCH_EN = RETURN_REG_EN;
  assign ALU_OUTREG_EN = RETURN_REG_EN;
  assign IR_LATCH_EN = NPC1_LATCH_EN;
  assign RegA_LATCH_EN = RD1;
  assign RegB_LATCH_EN = RD2;
  assign n209 = Rst;

  DFFS_X1 \cw1_reg[20]  ( .D(cw[6]), .CK(N442), .SN(n219), .Q(NPC1_LATCH_EN)
         );
  DFFR_X1 \cw1_reg[19]  ( .D(cw[19]), .CK(N442), .RN(n218), .Q(cw1[19]) );
  DFFR_X1 \cw1_reg[18]  ( .D(cw[18]), .CK(N442), .RN(n217), .Q(cw1[18]) );
  DFFR_X1 \cw1_reg[17]  ( .D(cw[17]), .CK(N442), .RN(n217), .Q(cw1[17]) );
  DFFR_X1 \cw1_reg[16]  ( .D(cw[5]), .CK(N442), .RN(n217), .Q(cw1[16]) );
  DFFR_X1 \cw1_reg[15]  ( .D(cw[15]), .CK(N442), .RN(n215), .Q(cw1[15]) );
  DFFR_X1 \cw1_reg[14]  ( .D(cw[14]), .CK(N442), .RN(n217), .Q(cw1[14]) );
  DFFR_X1 \cw1_reg[13]  ( .D(cw[7]), .CK(N442), .RN(n215), .Q(cw1[13]) );
  DFFR_X1 \cw1_reg[12]  ( .D(cw[5]), .CK(N442), .RN(n215), .Q(cw1[12]) );
  DFFR_X1 \cw1_reg[11]  ( .D(cw[15]), .CK(N442), .RN(n215), .Q(cw1[11]) );
  DFFR_X1 \cw1_reg[10]  ( .D(cw[8]), .CK(N442), .RN(n218), .Q(cw1[10]) );
  DFFR_X1 \cw1_reg[9]  ( .D(cw[9]), .CK(N442), .RN(n213), .Q(cw1[9]) );
  DFFR_X1 \cw1_reg[8]  ( .D(cw[8]), .CK(N442), .RN(n215), .Q(cw1[8]) );
  DFFR_X1 \cw1_reg[7]  ( .D(cw[7]), .CK(N442), .RN(n219), .Q(cw1[7]) );
  DFFR_X1 \cw1_reg[6]  ( .D(cw[6]), .CK(N442), .RN(n213), .Q(cw1[6]) );
  DFFR_X1 \cw1_reg[5]  ( .D(cw[5]), .CK(N442), .RN(n213), .Q(cw1[5]) );
  DFFR_X1 \cw1_reg[4]  ( .D(cw[4]), .CK(N442), .RN(n219), .Q(cw1[4]) );
  DFFR_X1 \cw1_reg[3]  ( .D(cw[8]), .CK(N442), .RN(n216), .Q(cw1[3]) );
  DFFR_X1 \cw1_reg[2]  ( .D(cw[2]), .CK(N442), .RN(n218), .Q(cw1[2]) );
  DFFR_X1 \cw1_reg[1]  ( .D(cw[9]), .CK(N442), .RN(n219), .Q(cw1[1]) );
  DFFR_X1 \cw1_reg[0]  ( .D(cw[2]), .CK(N442), .RN(n214), .Q(cw1[0]) );
  DFF_X1 \cw2_reg2[15]  ( .D(n161), .CK(Clk), .Q(cw2[15]) );
  DFF_X1 \cw2_reg2[14]  ( .D(n159), .CK(Clk), .Q(cw2[14]) );
  DFF_X1 \cw2_reg2[13]  ( .D(n157), .CK(Clk), .Q(cw2[13]) );
  DFF_X1 \cw2_reg2[12]  ( .D(n155), .CK(Clk), .Q(cw2[12]) );
  DFF_X1 \cw2_reg2[11]  ( .D(n153), .CK(Clk), .Q(cw2[11]) );
  DFF_X1 \cw2_reg2[10]  ( .D(n151), .CK(Clk), .Q(cw2[10]) );
  DFF_X1 \cw2_reg2[9]  ( .D(n149), .CK(Clk), .Q(cw2[9]) );
  DFF_X1 \cw2_reg2[8]  ( .D(n147), .CK(Clk), .Q(cw2[8]) );
  DFF_X1 \cw2_reg2[7]  ( .D(n145), .CK(Clk), .Q(cw2[7]) );
  DFF_X1 \cw2_reg2[6]  ( .D(n143), .CK(Clk), .Q(cw2[6]) );
  DFF_X1 \cw2_reg2[5]  ( .D(n141), .CK(Clk), .Q(cw2[5]) );
  DFF_X1 \cw2_reg2[4]  ( .D(n139), .CK(Clk), .Q(cw2[4]) );
  DFF_X1 \cw2_reg2[3]  ( .D(n137), .CK(Clk), .Q(cw2[3]) );
  DFF_X1 \cw2_reg2[2]  ( .D(n135), .CK(Clk), .Q(cw2[2]) );
  DFF_X1 \cw2_reg2[1]  ( .D(n133), .CK(Clk), .Q(cw2[1]) );
  DFF_X1 \cw2_reg2[0]  ( .D(n131), .CK(Clk), .Q(cw2[0]) );
  DFF_X1 \cw1_reg2[20]  ( .D(n129), .CK(Clk), .Q(NPC1_LATCH_EN) );
  DFF_X1 \cw1_reg2[19]  ( .D(n127), .CK(Clk), .Q(cw1[19]) );
  DFFR_X1 \cw2_reg[19]  ( .D(cw1[19]), .CK(N442), .RN(n219), .Q(RD1) );
  DFF_X1 \cw1_reg2[18]  ( .D(n124), .CK(Clk), .Q(cw1[18]) );
  DFFR_X1 \cw2_reg[18]  ( .D(cw1[18]), .CK(N442), .RN(n214), .Q(RD2) );
  DFF_X1 \cw1_reg2[17]  ( .D(n121), .CK(Clk), .Q(cw1[17]) );
  DFFR_X1 \cw2_reg[17]  ( .D(cw1[17]), .CK(N442), .RN(n213), .Q(
        RegIMM_LATCH_EN) );
  DFFR_X1 \cw2_reg[16]  ( .D(cw1[16]), .CK(N442), .RN(n214), .Q(Reg_RD1_EN) );
  DFFR_X1 \cw2_reg[15]  ( .D(cw1[15]), .CK(N442), .RN(n214), .Q(cw2[15]) );
  DFFR_X1 \cw2_reg[14]  ( .D(cw1[14]), .CK(N442), .RN(n214), .Q(cw2[14]) );
  DFF_X1 \cw1_reg2[12]  ( .D(n103), .CK(Clk), .Q(cw1[12]) );
  DFFR_X1 \cw2_reg[12]  ( .D(cw1[12]), .CK(N442), .RN(n217), .Q(cw2[12]) );
  DFFR_X1 \cw3_reg[12]  ( .D(cw2[12]), .CK(N442), .RN(n216), .Q(Reg_RD2_EN) );
  DFF_X1 \cw1_reg2[11]  ( .D(n99), .CK(Clk), .Q(cw1[11]) );
  DFFR_X1 \cw2_reg[11]  ( .D(cw1[11]), .CK(N442), .RN(n214), .Q(cw2[11]) );
  DFFR_X1 \cw3_reg[11]  ( .D(cw2[11]), .CK(N442), .RN(n215), .Q(JUMP_en) );
  DFF_X1 \cw1_reg2[10]  ( .D(n95), .CK(Clk), .Q(cw1[10]) );
  DFFR_X1 \cw2_reg[10]  ( .D(cw1[10]), .CK(N442), .RN(n214), .Q(cw2[10]) );
  DFFR_X1 \cw3_reg[10]  ( .D(cw2[10]), .CK(N442), .RN(n217), .Q(cw3[10]) );
  DFFR_X1 \cw4_reg[10]  ( .D(cw3[10]), .CK(N442), .RN(n218), .Q(DRAM_WE) );
  DFF_X1 \cw1_reg2[9]  ( .D(n90), .CK(Clk), .Q(cw1[9]) );
  DFFR_X1 \cw2_reg[9]  ( .D(cw1[9]), .CK(N442), .RN(n218), .Q(cw2[9]) );
  DFFR_X1 \cw3_reg[9]  ( .D(cw2[9]), .CK(N442), .RN(n217), .Q(cw3[9]) );
  DFF_X1 \cw1_reg2[8]  ( .D(n85), .CK(Clk), .Q(cw1[8]) );
  DFFR_X1 \cw2_reg[8]  ( .D(cw1[8]), .CK(N442), .RN(n218), .Q(cw2[8]) );
  DFFR_X1 \cw3_reg[8]  ( .D(cw2[8]), .CK(N442), .RN(n217), .Q(cw3[8]) );
  DFF_X1 \cw1_reg2[7]  ( .D(n80), .CK(Clk), .Q(cw1[7]) );
  DFFR_X1 \cw2_reg[7]  ( .D(cw1[7]), .CK(N442), .RN(n218), .Q(cw2[7]) );
  DFFR_X1 \cw3_reg[7]  ( .D(cw2[7]), .CK(N442), .RN(n218), .Q(cw3[7]) );
  DFF_X1 \cw1_reg2[6]  ( .D(n75), .CK(Clk), .Q(cw1[6]) );
  DFFR_X1 \cw2_reg[6]  ( .D(cw1[6]), .CK(N442), .RN(n217), .Q(cw2[6]) );
  DFFR_X1 \cw3_reg[6]  ( .D(cw2[6]), .CK(N442), .RN(n214), .Q(cw3[6]) );
  DFFR_X1 \cw4_reg[6]  ( .D(cw3[6]), .CK(N442), .RN(n218), .Q(PC_LATCH_EN) );
  DFF_X1 \cw1_reg2[5]  ( .D(n70), .CK(Clk), .Q(cw1[5]) );
  DFFR_X1 \cw2_reg[5]  ( .D(cw1[5]), .CK(N442), .RN(n217), .Q(cw2[5]) );
  DFFR_X1 \cw3_reg[5]  ( .D(cw2[5]), .CK(N442), .RN(n214), .Q(cw3[5]) );
  DFFR_X1 \cw4_reg[5]  ( .D(cw3[5]), .CK(N442), .RN(n214), .Q(Reg_RD3_EN) );
  DFF_X1 \cw1_reg2[4]  ( .D(n65), .CK(Clk), .Q(cw1[4]) );
  DFFR_X1 \cw2_reg[4]  ( .D(cw1[4]), .CK(N442), .RN(n213), .Q(cw2[4]) );
  DFFR_X1 \cw3_reg[4]  ( .D(cw2[4]), .CK(N442), .RN(n216), .Q(cw3[4]) );
  DFFR_X1 \cw4_reg[4]  ( .D(cw3[4]), .CK(N442), .RN(n214), .Q(
        write_stop_if_branch) );
  DFF_X1 \cw1_reg2[3]  ( .D(n60), .CK(Clk), .Q(cw1[3]) );
  DFFR_X1 \cw2_reg[3]  ( .D(cw1[3]), .CK(N442), .RN(n213), .Q(cw2[3]) );
  DFFR_X1 \cw3_reg[3]  ( .D(cw2[3]), .CK(N442), .RN(n216), .Q(cw3[3]) );
  DFFR_X1 \cw4_reg[3]  ( .D(cw3[3]), .CK(N442), .RN(n216), .Q(cw4[3]) );
  DFF_X1 \cw1_reg2[2]  ( .D(n54), .CK(Clk), .Q(cw1[2]) );
  DFFR_X1 \cw2_reg[2]  ( .D(cw1[2]), .CK(N442), .RN(n213), .Q(cw2[2]) );
  DFFR_X1 \cw3_reg[2]  ( .D(cw2[2]), .CK(N442), .RN(n215), .Q(cw3[2]) );
  DFFR_X1 \cw4_reg[2]  ( .D(cw3[2]), .CK(N442), .RN(n216), .Q(cw4[2]) );
  DFFR_X1 \cw5_reg[2]  ( .D(cw4[2]), .CK(N442), .RN(n213), .Q(RF_WE) );
  DFF_X1 \cw1_reg2[1]  ( .D(n48), .CK(Clk), .Q(cw1[1]) );
  DFFR_X1 \cw2_reg[1]  ( .D(cw1[1]), .CK(N442), .RN(n213), .Q(cw2[1]) );
  DFFR_X1 \cw3_reg[1]  ( .D(cw2[1]), .CK(N442), .RN(n216), .Q(cw3[1]) );
  DFFR_X1 \cw4_reg[1]  ( .D(cw3[1]), .CK(N442), .RN(n217), .Q(cw4[1]) );
  DFFR_X1 \cw5_reg[1]  ( .D(cw4[1]), .CK(N442), .RN(n213), .Q(WB_MUX_ADD_SEL)
         );
  DFF_X1 \cw1_reg2[0]  ( .D(n42), .CK(Clk), .Q(cw1[0]) );
  DFFR_X1 \cw2_reg[0]  ( .D(cw1[0]), .CK(N442), .RN(n213), .Q(cw2[0]) );
  DFFR_X1 \cw3_reg[0]  ( .D(cw2[0]), .CK(N442), .RN(n216), .Q(cw3[0]) );
  DFFR_X1 \cw4_reg[0]  ( .D(cw3[0]), .CK(N442), .RN(n216), .Q(cw4[0]) );
  DFFR_X1 \cw5_reg[0]  ( .D(cw4[0]), .CK(N442), .RN(n216), .Q(WR) );
  DFFR_X1 \cw2_reg[13]  ( .D(cw1[13]), .CK(N442), .RN(n215), .Q(cw2[13]) );
  DFFR_X1 \cw5_reg[3]  ( .D(cw4[3]), .CK(N442), .RN(n215), .Q(WB_MUX_SEL) );
  DFFR_X1 \cw4_reg[9]  ( .D(cw3[9]), .CK(N442), .RN(n218), .Q(ALU_OUT2_SEL) );
  DFFR_X1 \cw4_reg[8]  ( .D(cw3[8]), .CK(N442), .RN(n218), .Q(LMD_LATCH_EN) );
  DFFR_X1 \cw4_reg[7]  ( .D(cw3[7]), .CK(N442), .RN(n216), .Q(Alu_outreg2_en)
         );
  DFFR_X1 \cw3_reg[13]  ( .D(cw2[13]), .CK(N442), .RN(n215), .Q(RETURN_REG_EN)
         );
  DFFR_X1 \cw3_reg[14]  ( .D(cw2[14]), .CK(N442), .RN(n215), .Q(MUXB_SEL) );
  SDFFR_X1 \cw3_reg[15]  ( .D(1'b0), .SI(cw2[15]), .SE(1'b1), .CK(N442), .RN(
        n219), .Q(MUXA_SEL) );
  DFF_X1 \cw2_reg2[16]  ( .D(n163), .CK(Clk), .Q(Reg_RD1_EN) );
  DFF_X1 \cw1_reg2[16]  ( .D(n118), .CK(Clk), .Q(cw1[16]) );
  DFF_X1 \cw1_reg2[15]  ( .D(n115), .CK(Clk), .Q(cw1[15]) );
  DFF_X1 \cw1_reg2[14]  ( .D(n111), .CK(Clk), .Q(cw1[14]) );
  DFF_X1 \cw1_reg2[13]  ( .D(n107), .CK(Clk), .Q(cw1[13]) );
  DFF_X2 \cw2_reg2[18]  ( .D(n167), .CK(Clk), .Q(RD2) );
  DFF_X2 \cw2_reg2[19]  ( .D(n169), .CK(Clk), .Q(RD1) );
  DFF_X2 \cw2_reg2[17]  ( .D(n165), .CK(Clk), .Q(RegIMM_LATCH_EN) );
  INV_X2 U89 ( .A(Clk), .ZN(N442) );
  NAND3_X1 U90 ( .A1(IR_IN_26), .A2(n64), .A3(IR_IN_31), .ZN(n22) );
  OAI33_X1 U91 ( .A1(n28), .A2(IR_IN_27), .A3(n30), .B1(n58), .B2(IR_IN_29), 
        .B3(IR_IN_26), .ZN(n69) );
  NAND2_X1 U5 ( .A1(n25), .A2(n26), .ZN(cw[7]) );
  INV_X1 U6 ( .A(n26), .ZN(cw[5]) );
  OR2_X1 U7 ( .A1(cw[5]), .A2(cw[9]), .ZN(cw[2]) );
  INV_X1 U8 ( .A(n25), .ZN(cw[15]) );
  NOR2_X1 U9 ( .A1(flush), .A2(n20), .ZN(n165) );
  NOR2_X1 U10 ( .A1(flush), .A2(n21), .ZN(n163) );
  NAND2_X1 U11 ( .A1(n21), .A2(n20), .ZN(RegAluOpCodeGen_EN) );
  NOR2_X1 U12 ( .A1(n32), .A2(cw[18]), .ZN(n26) );
  NAND2_X1 U13 ( .A1(n31), .A2(n26), .ZN(cw[19]) );
  NAND2_X1 U14 ( .A1(n64), .A2(n29), .ZN(n25) );
  NOR2_X1 U15 ( .A1(n30), .A2(n25), .ZN(cw[9]) );
  INV_X1 U16 ( .A(n22), .ZN(cw[8]) );
  OR2_X1 U17 ( .A1(n32), .A2(cw[15]), .ZN(cw[14]) );
  OR2_X1 U18 ( .A1(n32), .A2(cw[4]), .ZN(cw[17]) );
  BUF_X1 U19 ( .A(n209), .Z(n211) );
  BUF_X1 U20 ( .A(n209), .Z(n212) );
  AND2_X1 U21 ( .A1(RD1), .A2(n220), .ZN(n169) );
  AND2_X1 U22 ( .A1(RD2), .A2(n221), .ZN(n167) );
  AND2_X1 U23 ( .A1(NPC1_LATCH_EN), .A2(n220), .ZN(n129) );
  AND2_X1 U24 ( .A1(cw1[13]), .A2(n220), .ZN(n107) );
  AND2_X1 U25 ( .A1(cw1[14]), .A2(n220), .ZN(n111) );
  AND2_X1 U26 ( .A1(cw1[15]), .A2(n220), .ZN(n115) );
  AND2_X1 U27 ( .A1(cw1[16]), .A2(n220), .ZN(n118) );
  AND2_X1 U28 ( .A1(cw1[0]), .A2(n220), .ZN(n42) );
  AND2_X1 U29 ( .A1(cw1[1]), .A2(n221), .ZN(n48) );
  AND2_X1 U30 ( .A1(cw1[2]), .A2(n221), .ZN(n54) );
  AND2_X1 U31 ( .A1(cw1[3]), .A2(n220), .ZN(n60) );
  AND2_X1 U32 ( .A1(cw1[4]), .A2(n221), .ZN(n65) );
  AND2_X1 U33 ( .A1(cw1[5]), .A2(n220), .ZN(n70) );
  AND2_X1 U34 ( .A1(cw1[12]), .A2(n220), .ZN(n103) );
  AND2_X1 U35 ( .A1(cw1[17]), .A2(n220), .ZN(n121) );
  AND2_X1 U36 ( .A1(cw1[18]), .A2(n220), .ZN(n124) );
  AND2_X1 U37 ( .A1(cw1[19]), .A2(n220), .ZN(n127) );
  AND2_X1 U38 ( .A1(cw2[0]), .A2(n220), .ZN(n131) );
  AND2_X1 U39 ( .A1(cw2[1]), .A2(n220), .ZN(n133) );
  AND2_X1 U40 ( .A1(cw2[2]), .A2(n221), .ZN(n135) );
  AND2_X1 U41 ( .A1(cw2[3]), .A2(n221), .ZN(n137) );
  AND2_X1 U42 ( .A1(cw2[4]), .A2(n221), .ZN(n139) );
  AND2_X1 U43 ( .A1(cw2[5]), .A2(n221), .ZN(n141) );
  AND2_X1 U44 ( .A1(cw2[6]), .A2(n221), .ZN(n143) );
  AND2_X1 U45 ( .A1(cw2[7]), .A2(n221), .ZN(n145) );
  AND2_X1 U46 ( .A1(cw2[8]), .A2(n221), .ZN(n147) );
  AND2_X1 U47 ( .A1(cw2[9]), .A2(n221), .ZN(n149) );
  AND2_X1 U48 ( .A1(cw2[10]), .A2(n221), .ZN(n151) );
  AND2_X1 U49 ( .A1(cw2[11]), .A2(n221), .ZN(n153) );
  AND2_X1 U50 ( .A1(cw2[12]), .A2(n221), .ZN(n155) );
  AND2_X1 U51 ( .A1(cw2[13]), .A2(n220), .ZN(n157) );
  AND2_X1 U52 ( .A1(cw2[14]), .A2(n221), .ZN(n159) );
  AND2_X1 U53 ( .A1(cw2[15]), .A2(n221), .ZN(n161) );
  AND2_X1 U54 ( .A1(cw1[6]), .A2(n220), .ZN(n75) );
  AND2_X1 U55 ( .A1(cw1[7]), .A2(n220), .ZN(n80) );
  AND2_X1 U56 ( .A1(cw1[8]), .A2(n221), .ZN(n85) );
  AND2_X1 U57 ( .A1(cw1[9]), .A2(n220), .ZN(n90) );
  AND2_X1 U58 ( .A1(cw1[10]), .A2(n221), .ZN(n95) );
  AND2_X1 U59 ( .A1(cw1[11]), .A2(n221), .ZN(n99) );
  INV_X1 U60 ( .A(RegIMM_LATCH_EN), .ZN(n20) );
  INV_X1 U61 ( .A(Reg_RD1_EN), .ZN(n21) );
  NOR4_X1 U62 ( .A1(n41), .A2(n46), .A3(IR_IN[1]), .A4(n47), .ZN(n35) );
  INV_X1 U63 ( .A(IR_IN[0]), .ZN(n41) );
  INV_X1 U64 ( .A(IR_IN[5]), .ZN(n46) );
  NOR4_X1 U65 ( .A1(n27), .A2(IR_IN_28), .A3(IR_IN_29), .A4(IR_IN_30), .ZN(n64) );
  OAI221_X1 U66 ( .B1(IR_IN_31), .B2(n68), .C1(n28), .C2(n31), .A(n22), .ZN(
        n32) );
  AOI21_X1 U67 ( .B1(IR_IN_30), .B2(n69), .A(n73), .ZN(n68) );
  NOR3_X1 U68 ( .A1(n28), .A2(IR_IN_30), .A3(IR_IN_26), .ZN(n73) );
  NOR3_X1 U69 ( .A1(IR_IN_30), .A2(IR_IN_31), .A3(IR_IN_27), .ZN(n63) );
  NOR3_X1 U70 ( .A1(IR_IN[0]), .A2(IR_IN[3]), .A3(n47), .ZN(n34) );
  INV_X1 U71 ( .A(IR_IN_29), .ZN(n28) );
  NOR2_X1 U72 ( .A1(IR_IN[9]), .A2(IR_IN[8]), .ZN(n59) );
  OR4_X1 U73 ( .A1(IR_IN[10]), .A2(n52), .A3(n53), .A4(n55), .ZN(n47) );
  OR3_X1 U74 ( .A1(IR_IN[7]), .A2(IR_IN[6]), .A3(IR_IN[4]), .ZN(n53) );
  INV_X1 U75 ( .A(n63), .ZN(n52) );
  NAND4_X1 U76 ( .A1(n58), .A2(n28), .A3(n30), .A4(n59), .ZN(n55) );
  INV_X1 U77 ( .A(IR_IN_26), .ZN(n30) );
  INV_X1 U78 ( .A(n33), .ZN(cw[18]) );
  AOI221_X1 U79 ( .B1(IR_IN[5]), .B2(n34), .C1(n35), .C2(IR_IN[3]), .A(n36), 
        .ZN(n33) );
  INV_X1 U80 ( .A(n40), .ZN(n36) );
  OAI21_X1 U81 ( .B1(n34), .B2(n35), .A(IR_IN[2]), .ZN(n40) );
  INV_X1 U82 ( .A(IR_IN_27), .ZN(n27) );
  NAND2_X1 U83 ( .A1(n23), .A2(n24), .ZN(cw[6]) );
  NAND4_X1 U84 ( .A1(IR_IN_28), .A2(n27), .A3(n28), .A4(n29), .ZN(n23) );
  INV_X1 U85 ( .A(cw[7]), .ZN(n24) );
  INV_X1 U86 ( .A(IR_IN_28), .ZN(n58) );
  OAI21_X1 U87 ( .B1(IR_IN_29), .B2(n31), .A(n25), .ZN(cw[4]) );
  NAND2_X1 U88 ( .A1(IR_IN_28), .A2(n63), .ZN(n31) );
  INV_X1 U92 ( .A(IR_IN_31), .ZN(n29) );
  CLKBUF_X1 U93 ( .A(n211), .Z(n213) );
  CLKBUF_X1 U94 ( .A(n211), .Z(n214) );
  CLKBUF_X1 U95 ( .A(n211), .Z(n215) );
  CLKBUF_X1 U96 ( .A(n211), .Z(n216) );
  CLKBUF_X1 U97 ( .A(n212), .Z(n217) );
  CLKBUF_X1 U98 ( .A(n212), .Z(n218) );
  CLKBUF_X1 U99 ( .A(n212), .Z(n219) );
  INV_X1 U100 ( .A(flush), .ZN(n220) );
  INV_X1 U101 ( .A(flush), .ZN(n221) );
endmodule


module mux21_N32_0 ( A, B, SEL, Y );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Y;
  input SEL;
  wire   n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130;

  BUF_X1 U1 ( .A(n121), .Z(n130) );
  INV_X1 U2 ( .A(n130), .ZN(n118) );
  INV_X1 U3 ( .A(n130), .ZN(n117) );
  CLKBUF_X1 U4 ( .A(n121), .Z(n128) );
  BUF_X1 U5 ( .A(n119), .Z(n123) );
  CLKBUF_X1 U6 ( .A(n119), .Z(n122) );
  CLKBUF_X1 U7 ( .A(n119), .Z(n124) );
  BUF_X1 U8 ( .A(n120), .Z(n125) );
  CLKBUF_X1 U9 ( .A(n120), .Z(n127) );
  CLKBUF_X1 U10 ( .A(n120), .Z(n126) );
  CLKBUF_X1 U11 ( .A(n121), .Z(n129) );
  BUF_X1 U12 ( .A(SEL), .Z(n121) );
  CLKBUF_X1 U13 ( .A(SEL), .Z(n119) );
  CLKBUF_X1 U14 ( .A(SEL), .Z(n120) );
  INV_X1 U15 ( .A(n53), .ZN(Y[21]) );
  AOI22_X1 U16 ( .A1(A[21]), .A2(n117), .B1(B[21]), .B2(n126), .ZN(n53) );
  INV_X1 U17 ( .A(n43), .ZN(Y[30]) );
  AOI22_X1 U18 ( .A1(A[30]), .A2(n118), .B1(B[30]), .B2(n126), .ZN(n43) );
  INV_X1 U19 ( .A(n45), .ZN(Y[29]) );
  AOI22_X1 U20 ( .A1(A[29]), .A2(n118), .B1(B[29]), .B2(n124), .ZN(n45) );
  INV_X1 U21 ( .A(n46), .ZN(Y[28]) );
  AOI22_X1 U22 ( .A1(A[28]), .A2(n117), .B1(B[28]), .B2(n124), .ZN(n46) );
  INV_X1 U23 ( .A(n47), .ZN(Y[27]) );
  AOI22_X1 U24 ( .A1(A[27]), .A2(n117), .B1(B[27]), .B2(n124), .ZN(n47) );
  INV_X1 U25 ( .A(n48), .ZN(Y[26]) );
  AOI22_X1 U26 ( .A1(A[26]), .A2(n118), .B1(B[26]), .B2(n124), .ZN(n48) );
  INV_X1 U27 ( .A(n49), .ZN(Y[25]) );
  AOI22_X1 U28 ( .A1(A[25]), .A2(n117), .B1(B[25]), .B2(n125), .ZN(n49) );
  INV_X1 U29 ( .A(n50), .ZN(Y[24]) );
  AOI22_X1 U30 ( .A1(A[24]), .A2(n117), .B1(B[24]), .B2(n125), .ZN(n50) );
  INV_X1 U31 ( .A(n51), .ZN(Y[23]) );
  AOI22_X1 U32 ( .A1(A[23]), .A2(n118), .B1(B[23]), .B2(n125), .ZN(n51) );
  INV_X1 U33 ( .A(n52), .ZN(Y[22]) );
  AOI22_X1 U34 ( .A1(A[22]), .A2(n118), .B1(B[22]), .B2(n125), .ZN(n52) );
  INV_X1 U35 ( .A(n54), .ZN(Y[20]) );
  AOI22_X1 U36 ( .A1(A[20]), .A2(n118), .B1(B[20]), .B2(n126), .ZN(n54) );
  INV_X1 U37 ( .A(n56), .ZN(Y[19]) );
  AOI22_X1 U38 ( .A1(A[19]), .A2(n118), .B1(B[19]), .B2(n127), .ZN(n56) );
  INV_X1 U39 ( .A(n57), .ZN(Y[18]) );
  AOI22_X1 U40 ( .A1(A[18]), .A2(n117), .B1(B[18]), .B2(n127), .ZN(n57) );
  INV_X1 U41 ( .A(n58), .ZN(Y[17]) );
  AOI22_X1 U42 ( .A1(A[17]), .A2(n118), .B1(B[17]), .B2(n127), .ZN(n58) );
  INV_X1 U43 ( .A(n59), .ZN(Y[16]) );
  AOI22_X1 U44 ( .A1(A[16]), .A2(n117), .B1(B[16]), .B2(n127), .ZN(n59) );
  INV_X1 U45 ( .A(n60), .ZN(Y[15]) );
  AOI22_X1 U46 ( .A1(A[15]), .A2(n118), .B1(B[15]), .B2(n128), .ZN(n60) );
  INV_X1 U47 ( .A(n61), .ZN(Y[14]) );
  AOI22_X1 U48 ( .A1(A[14]), .A2(n117), .B1(B[14]), .B2(n128), .ZN(n61) );
  INV_X1 U49 ( .A(n62), .ZN(Y[13]) );
  AOI22_X1 U50 ( .A1(A[13]), .A2(n117), .B1(B[13]), .B2(n128), .ZN(n62) );
  INV_X1 U51 ( .A(n63), .ZN(Y[12]) );
  AOI22_X1 U52 ( .A1(A[12]), .A2(n118), .B1(B[12]), .B2(n128), .ZN(n63) );
  INV_X1 U53 ( .A(n64), .ZN(Y[11]) );
  AOI22_X1 U54 ( .A1(A[11]), .A2(n117), .B1(B[11]), .B2(n129), .ZN(n64) );
  INV_X1 U55 ( .A(n65), .ZN(Y[10]) );
  AOI22_X1 U56 ( .A1(A[10]), .A2(n117), .B1(B[10]), .B2(n129), .ZN(n65) );
  INV_X1 U57 ( .A(n66), .ZN(Y[0]) );
  AOI22_X1 U58 ( .A1(A[0]), .A2(n117), .B1(B[0]), .B2(n129), .ZN(n66) );
  INV_X1 U59 ( .A(n44), .ZN(Y[2]) );
  AOI22_X1 U60 ( .A1(A[2]), .A2(n118), .B1(B[2]), .B2(n123), .ZN(n44) );
  INV_X1 U61 ( .A(n55), .ZN(Y[1]) );
  AOI22_X1 U62 ( .A1(A[1]), .A2(n118), .B1(B[1]), .B2(n126), .ZN(n55) );
  INV_X1 U63 ( .A(n41), .ZN(Y[3]) );
  AOI22_X1 U64 ( .A1(A[3]), .A2(n118), .B1(B[3]), .B2(n123), .ZN(n41) );
  INV_X1 U65 ( .A(n37), .ZN(Y[7]) );
  AOI22_X1 U66 ( .A1(A[7]), .A2(n118), .B1(B[7]), .B2(n122), .ZN(n37) );
  INV_X1 U67 ( .A(n34), .ZN(Y[9]) );
  AOI22_X1 U68 ( .A1(A[9]), .A2(n118), .B1(n129), .B2(B[9]), .ZN(n34) );
  INV_X1 U69 ( .A(n40), .ZN(Y[4]) );
  AOI22_X1 U70 ( .A1(A[4]), .A2(n117), .B1(B[4]), .B2(n123), .ZN(n40) );
  INV_X1 U71 ( .A(n36), .ZN(Y[8]) );
  AOI22_X1 U72 ( .A1(A[8]), .A2(n117), .B1(B[8]), .B2(n122), .ZN(n36) );
  INV_X1 U73 ( .A(n38), .ZN(Y[6]) );
  AOI22_X1 U74 ( .A1(A[6]), .A2(n117), .B1(B[6]), .B2(n122), .ZN(n38) );
  INV_X1 U75 ( .A(n39), .ZN(Y[5]) );
  AOI22_X1 U76 ( .A1(A[5]), .A2(n118), .B1(B[5]), .B2(n122), .ZN(n39) );
  INV_X1 U77 ( .A(n42), .ZN(Y[31]) );
  AOI22_X1 U78 ( .A1(A[31]), .A2(n117), .B1(B[31]), .B2(n123), .ZN(n42) );
endmodule


module datapath_reg_size32 ( clk, rst, flush, RF1, RF2, WF1, EN_regA, EN_regB, 
        EN_regIMM, EN_regALUOP, EN_regRD1, EN_regNPC2, S1, S2, EN_regRET, 
        EN_regOUTALU, EN_regB2, EN_regRD2, EN_regALU2, EN_regLMD, EN_regRD3, 
        Sel_ret_alu, Sel_alu_lmd, sel_31_rd, NPC, IR_dp, OUT_DP, comp_branch_i, 
        immediate_branch, ADD_mem, DIN_mem, DOUT_mem );
  input [31:0] NPC;
  input [31:0] IR_dp;
  output [31:0] OUT_DP;
  output [31:0] immediate_branch;
  output [31:0] ADD_mem;
  output [31:0] DIN_mem;
  input [31:0] DOUT_mem;
  input clk, rst, flush, RF1, RF2, WF1, EN_regA, EN_regB, EN_regIMM,
         EN_regALUOP, EN_regRD1, EN_regNPC2, S1, S2, EN_regRET, EN_regOUTALU,
         EN_regB2, EN_regRD2, EN_regALU2, EN_regLMD, EN_regRD3, Sel_ret_alu,
         Sel_alu_lmd, sel_31_rd;
  output comp_branch_i;
  wire   jump_op, N40, N47, N49, N51, N53, N55, N56, add_sub_i, n1, n29, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n31, n32;
  wire   [4:0] add_w_rf;
  wire   [31:0] alu2_lmd;
  wire   [31:0] A;
  wire   [31:0] B;
  wire   [31:0] ext;
  wire   [31:0] out_A;
  wire   [31:0] out_b;
  wire   [31:0] npc2;
  wire   [16:0] aluopcode_reg_out;
  wire   [4:0] signal_rd_in;
  wire   [4:0] out_rd1;
  wire   [31:0] out_mux_1;
  wire   [31:0] out_mux_2;
  wire   [2:0] aluopcode_i;
  wire   [3:0] compare_code_i;
  wire   [2:0] shiftopcode_i;
  wire   [31:0] reg_alu_in;
  wire   [31:0] return_alu;
  wire   [4:0] out_rd2;
  wire   [31:0] return_out;
  wire   [31:0] out_ret_alu;
  wire   [31:0] alu2;
  wire   [31:0] lmd;
  wire   [4:0] rd3;
  tri   RF1;
  tri   RF2;
  tri   EN_regA;
  tri   EN_regB;
  tri   EN_regIMM;
  tri   EN_regRD1;
  assign OUT_DP[31] = ADD_mem[31];
  assign OUT_DP[30] = ADD_mem[30];
  assign OUT_DP[29] = ADD_mem[29];
  assign OUT_DP[28] = ADD_mem[28];
  assign OUT_DP[27] = ADD_mem[27];
  assign OUT_DP[26] = ADD_mem[26];
  assign OUT_DP[25] = ADD_mem[25];
  assign OUT_DP[24] = ADD_mem[24];
  assign OUT_DP[23] = ADD_mem[23];
  assign OUT_DP[22] = ADD_mem[22];
  assign OUT_DP[21] = ADD_mem[21];
  assign OUT_DP[20] = ADD_mem[20];
  assign OUT_DP[19] = ADD_mem[19];
  assign OUT_DP[18] = ADD_mem[18];
  assign OUT_DP[17] = ADD_mem[17];
  assign OUT_DP[16] = ADD_mem[16];
  assign OUT_DP[15] = ADD_mem[15];
  assign OUT_DP[14] = ADD_mem[14];
  assign OUT_DP[13] = ADD_mem[13];
  assign OUT_DP[12] = ADD_mem[12];
  assign OUT_DP[11] = ADD_mem[11];
  assign OUT_DP[10] = ADD_mem[10];
  assign OUT_DP[9] = ADD_mem[9];
  assign OUT_DP[8] = ADD_mem[8];
  assign OUT_DP[7] = ADD_mem[7];
  assign OUT_DP[6] = ADD_mem[6];
  assign OUT_DP[5] = ADD_mem[5];
  assign OUT_DP[4] = ADD_mem[4];
  assign OUT_DP[3] = ADD_mem[3];
  assign OUT_DP[2] = ADD_mem[2];
  assign OUT_DP[1] = ADD_mem[1];
  assign OUT_DP[0] = ADD_mem[0];
  assign n29 = rst;

  DLH_X1 jump_op_reg ( .G(N56), .D(N40), .Q(jump_op) );
  DLL_X1 \signal_rd_in_reg[4]  ( .D(N55), .GN(N56), .Q(signal_rd_in[4]) );
  DLL_X1 \signal_rd_in_reg[3]  ( .D(N53), .GN(N56), .Q(signal_rd_in[3]) );
  DLL_X1 \signal_rd_in_reg[2]  ( .D(N51), .GN(N56), .Q(signal_rd_in[2]) );
  DLL_X1 \signal_rd_in_reg[1]  ( .D(N49), .GN(N56), .Q(signal_rd_in[1]) );
  DLL_X1 \signal_rd_in_reg[0]  ( .D(N47), .GN(N56), .Q(signal_rd_in[0]) );
  NOR4_X2 U18 ( .A1(IR_dp[26]), .A2(n24), .A3(IR_dp[28]), .A4(IR_dp[27]), .ZN(
        n19) );
  NAND3_X1 U23 ( .A1(n15), .A2(n16), .A3(IR_dp[28]), .ZN(n14) );
  register_file_NBIT32_row32 rf ( .CLK(clk), .RESET(n31), .ENABLE(1'b1), .RD1(
        RF1), .RD2(RF2), .WR(WF1), .ADD_WR(add_w_rf), .ADD_RD1(IR_dp[25:21]), 
        .ADD_RD2(IR_dp[20:16]), .DATAIN(alu2_lmd), .OUT1(A), .OUT2(B) );
  SIG_EXT_BITS32 estensione_segno ( .EXT_UNSIGNED(1'b1), .EXT_FOR_J(jump_op), 
        .S_IN(IR_dp), .S_OUT(ext) );
  registro_N32_0 reg_A ( .data(A), .enable(EN_regA), .clock(clk), .clear(n1), 
        .Q(out_A) );
  registro_N32_8 reg_B ( .data(B), .enable(EN_regB), .clock(clk), .clear(n1), 
        .Q(out_b) );
  registro_N32_7 reg_NPC2 ( .data(NPC), .enable(EN_regNPC2), .clock(clk), 
        .clear(n31), .Q(npc2) );
  registro_N32_6 reg_IMMEDIATE ( .data(ext), .enable(EN_regIMM), .clock(clk), 
        .clear(n31), .Q(immediate_branch) );
  registro_N17 reg_aluopcode ( .data({IR_dp[31:26], IR_dp[10:0]}), .enable(
        EN_regALUOP), .clock(clk), .clear(n31), .Q(aluopcode_reg_out) );
  registro_N5_0 reg_rd1 ( .data(signal_rd_in), .enable(EN_regRD1), .clock(clk), 
        .clear(n1), .Q(out_rd1) );
  mux21_N32_4 mux_in1_A ( .A(out_A), .B(npc2), .SEL(S1), .Y(out_mux_1) );
  mux21_N32_3 mux_in1_B ( .A(out_b), .B(immediate_branch), .SEL(S2), .Y(
        out_mux_2) );
  ALU_N32 alu_dlx ( .AluOpCode(aluopcode_i), .CompareOpCode(compare_code_i), 
        .Add_subn(add_sub_i), .ShiftOpCode(shiftopcode_i), .DATA1(out_mux_1), 
        .DATA2(out_mux_2), .OUTALU(reg_alu_in), .return_address(return_alu), 
        .CompBranch(comp_branch_i) );
  AluOpCodeGen alu_opcode_generator ( .IR_opcode(aluopcode_reg_out[16:11]), 
        .IR_func(aluopcode_reg_out[10:0]), .AluOpCode(aluopcode_i), .Add_Subn(
        add_sub_i), .CompareCode(compare_code_i), .ShiftOpCode(shiftopcode_i)
         );
  registro_N32_5 reg_alu_out ( .data(reg_alu_in), .enable(EN_regOUTALU), 
        .clock(clk), .clear(n31), .Q(ADD_mem) );
  registro_N32_4 reg_b2 ( .data(out_b), .enable(EN_regB2), .clock(clk), 
        .clear(n31), .Q(DIN_mem) );
  registro_N5_2 reg_rd2 ( .data(out_rd1), .enable(EN_regRD2), .clock(clk), 
        .clear(n31), .Q(out_rd2) );
  registro_N32_3 reg_return ( .data(return_alu), .enable(EN_regRET), .clock(
        clk), .clear(n31), .Q(return_out) );
  mux21_N32_2 mux_ret_alu ( .A(ADD_mem), .B(return_out), .SEL(Sel_ret_alu), 
        .Y(out_ret_alu) );
  registro_N32_2 reg_alu2 ( .data(out_ret_alu), .enable(EN_regALU2), .clock(
        clk), .clear(n31), .Q(alu2) );
  registro_N32_1 reg_lmd ( .data(DOUT_mem), .enable(EN_regLMD), .clock(clk), 
        .clear(n31), .Q(lmd) );
  registro_N5_1 reg_rd3 ( .data(out_rd2), .enable(EN_regRD3), .clock(clk), 
        .clear(n31), .Q(rd3) );
  mux21_N32_1 mux_lmd_alu ( .A(alu2), .B(lmd), .SEL(Sel_alu_lmd), .Y(alu2_lmd)
         );
  mux21_N5 mux_address_write ( .A(rd3), .B({1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), 
        .SEL(sel_31_rd), .Y(add_w_rf) );
  NOR2_X1 U3 ( .A1(flush), .A2(n32), .ZN(n1) );
  INV_X2 U4 ( .A(n32), .ZN(n31) );
  INV_X1 U5 ( .A(n19), .ZN(n18) );
  INV_X1 U6 ( .A(n29), .ZN(n32) );
  INV_X1 U7 ( .A(n15), .ZN(n24) );
  NOR3_X1 U8 ( .A1(IR_dp[31]), .A2(IR_dp[30]), .A3(IR_dp[29]), .ZN(n15) );
  NOR3_X1 U9 ( .A1(n24), .A2(IR_dp[28]), .A3(n16), .ZN(N40) );
  NAND2_X1 U10 ( .A1(n13), .A2(n14), .ZN(N56) );
  INV_X1 U11 ( .A(N40), .ZN(n13) );
  INV_X1 U12 ( .A(IR_dp[27]), .ZN(n16) );
  INV_X1 U13 ( .A(n23), .ZN(N47) );
  AOI22_X1 U14 ( .A1(IR_dp[16]), .A2(n18), .B1(IR_dp[11]), .B2(n19), .ZN(n23)
         );
  INV_X1 U15 ( .A(n22), .ZN(N49) );
  AOI22_X1 U16 ( .A1(IR_dp[17]), .A2(n18), .B1(IR_dp[12]), .B2(n19), .ZN(n22)
         );
  INV_X1 U17 ( .A(n21), .ZN(N51) );
  AOI22_X1 U19 ( .A1(IR_dp[18]), .A2(n18), .B1(IR_dp[13]), .B2(n19), .ZN(n21)
         );
  INV_X1 U20 ( .A(n20), .ZN(N53) );
  AOI22_X1 U21 ( .A1(IR_dp[19]), .A2(n18), .B1(IR_dp[14]), .B2(n19), .ZN(n20)
         );
  INV_X1 U22 ( .A(n17), .ZN(N55) );
  AOI22_X1 U24 ( .A1(IR_dp[20]), .A2(n18), .B1(IR_dp[15]), .B2(n19), .ZN(n17)
         );
endmodule


module DLX_IR_SIZE32_PC_SIZE32 ( Clk, Rst, dram_RD, dram_WR, dram_ADD, 
        dram_DIN, dram_DOUT, iram_Addr, iram_Dout );
  output [31:0] dram_ADD;
  output [31:0] dram_DIN;
  input [31:0] dram_DOUT;
  output [31:0] iram_Addr;
  input [31:0] iram_Dout;
  input Clk, Rst;
  output dram_RD, dram_WR;
  wire   wr_i, MUXA_SEL_i, MUXB_SEL_i, RETURN_REG_EN_i, ALU_OUTREG_EN_i,
         B2_EN_i, en_RD2_i, Alu_outreg2_en_i, LMD_LATCH_EN_i, en_RD3_i,
         sel_alu_ret_i, WB_MUX_SEL_i, wb_mux_add_sel_i, comp_branch_dp,
         JUMP_EN_i, wr_cu, write_stop_if_branch_i, net3527, net3526, net3525,
         net3524, net3523, net3522, net3521, net3520, net3519, net3518,
         net3517, net3516, net3515, net3514, net3513, net3512, net3511,
         net3510, net3509, net3508, net3507, net3506, net3505, net3504,
         net3503, net3502, net3501, net3500, net3499, net3498, net3497,
         net3496, net3495, net3494, net3493, net3492, net3491, net3490,
         net3489, net3488, net3487, net3486, net3485, net3484, net3483,
         net3482, net3481, net3480, net3479, net3478, net3477, net3476,
         net3475, net3474, net3473, net3472, net3471, net3470, net3469,
         net3468, net3467, net3466, net3465, net3464, net3431, net3430,
         net3429, net3428, net3427, net3426, net3425, net3424, net3423,
         net3422, net3421, net3420, net3419, net3418, net3417, net3416,
         net3415, net3414, net3413, net3412, net3411, net3410, net3409,
         net3408, net3407, net3406, net3405, net3404, net3403, net3402,
         net3401, net3400, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n1225,
         n1230, n1233, n1238, n1244, n1284, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435;
  wire   [31:0] out_NPC;
  wire   [31:0] IR;
  wire   [31:0] immediate;
  wire   [31:0] PC;
  wire   [31:0] PC_BUS;
  wire   [31:0] in_NPC;
  wire   [31:0] npc2;
  wire   [31:0] pc_jump;
  tri   en_RD1_i;
wand  rd1_i;
wand  rd2_i;
wand  RegA_LATCH_EN_i;
wand  RegB_LATCH_EN_i;
wand  RegIMM_LATCH_EN_i;
wand  NPC1_LATCH_EN_i;
  assign n1244 = Rst;

  DFFR_X1 \npc2_reg[0]  ( .D(n296), .CK(Clk), .RN(n1422), .Q(npc2[0]), .QN(
        net3400) );
  DFFR_X1 \npc2_reg[31]  ( .D(n293), .CK(Clk), .RN(n1422), .Q(npc2[31]), .QN(
        net3431) );
  DFFR_X1 \npc2_reg[1]  ( .D(n290), .CK(Clk), .RN(n1418), .Q(npc2[1]), .QN(
        net3401) );
  DFFR_X1 \npc2_reg[2]  ( .D(n288), .CK(Clk), .RN(n1418), .Q(npc2[2]), .QN(
        net3402) );
  DFFR_X1 \npc2_reg[3]  ( .D(n286), .CK(Clk), .RN(n1418), .Q(npc2[3]), .QN(
        net3403) );
  DFFR_X1 \npc2_reg[4]  ( .D(n284), .CK(Clk), .RN(n1419), .Q(npc2[4]), .QN(
        net3404) );
  DFFR_X1 \npc2_reg[5]  ( .D(n282), .CK(Clk), .RN(n1420), .Q(npc2[5]), .QN(
        net3405) );
  DFFR_X1 \npc2_reg[6]  ( .D(n280), .CK(Clk), .RN(n1419), .Q(npc2[6]), .QN(
        net3406) );
  DFFR_X1 \npc2_reg[7]  ( .D(n278), .CK(Clk), .RN(n1418), .Q(npc2[7]), .QN(
        net3407) );
  DFFR_X1 \npc2_reg[8]  ( .D(n276), .CK(Clk), .RN(n1418), .Q(npc2[8]), .QN(
        net3408) );
  DFFR_X1 \npc2_reg[9]  ( .D(n274), .CK(Clk), .RN(n1419), .Q(npc2[9]), .QN(
        net3409) );
  DFFR_X1 \npc2_reg[10]  ( .D(n272), .CK(Clk), .RN(n1418), .Q(npc2[10]), .QN(
        net3410) );
  DFFR_X1 \npc2_reg[11]  ( .D(n270), .CK(Clk), .RN(n1418), .Q(npc2[11]), .QN(
        net3411) );
  DFFR_X1 \npc2_reg[12]  ( .D(n268), .CK(Clk), .RN(n1419), .Q(npc2[12]), .QN(
        net3412) );
  DFFR_X1 \npc2_reg[13]  ( .D(n266), .CK(Clk), .RN(n1419), .Q(npc2[13]), .QN(
        net3413) );
  DFFR_X1 \npc2_reg[14]  ( .D(n264), .CK(Clk), .RN(n1419), .Q(npc2[14]), .QN(
        net3414) );
  DFFR_X1 \npc2_reg[15]  ( .D(n262), .CK(Clk), .RN(n1419), .Q(npc2[15]), .QN(
        net3415) );
  DFFR_X1 \npc2_reg[16]  ( .D(n260), .CK(Clk), .RN(n1420), .Q(npc2[16]), .QN(
        net3416) );
  DFFR_X1 \npc2_reg[17]  ( .D(n258), .CK(Clk), .RN(n1420), .Q(npc2[17]), .QN(
        net3417) );
  DFFR_X1 \npc2_reg[18]  ( .D(n256), .CK(Clk), .RN(n1423), .Q(npc2[18]), .QN(
        net3418) );
  DFFR_X1 \npc2_reg[19]  ( .D(n254), .CK(Clk), .RN(n1422), .Q(npc2[19]), .QN(
        net3419) );
  DFFR_X1 \npc2_reg[20]  ( .D(n252), .CK(Clk), .RN(n1422), .Q(npc2[20]), .QN(
        net3420) );
  DFFR_X1 \npc2_reg[21]  ( .D(n250), .CK(Clk), .RN(n1422), .Q(npc2[21]), .QN(
        net3421) );
  DFFR_X1 \npc2_reg[22]  ( .D(n248), .CK(Clk), .RN(n1418), .Q(npc2[22]), .QN(
        net3422) );
  DFFR_X1 \npc2_reg[23]  ( .D(n246), .CK(Clk), .RN(n1422), .Q(npc2[23]), .QN(
        net3423) );
  DFFR_X1 \npc2_reg[24]  ( .D(n244), .CK(Clk), .RN(n1422), .Q(npc2[24]), .QN(
        net3424) );
  DFFR_X1 \npc2_reg[25]  ( .D(n242), .CK(Clk), .RN(n1422), .Q(npc2[25]), .QN(
        net3425) );
  DFFR_X1 \npc2_reg[26]  ( .D(n240), .CK(Clk), .RN(n1419), .Q(npc2[26]), .QN(
        net3426) );
  DFFR_X1 \npc2_reg[27]  ( .D(n238), .CK(Clk), .RN(n1419), .Q(npc2[27]), .QN(
        net3427) );
  DFFR_X1 \npc2_reg[28]  ( .D(n236), .CK(Clk), .RN(n1422), .Q(npc2[28]), .QN(
        net3428) );
  DFFR_X1 \npc2_reg[29]  ( .D(n234), .CK(Clk), .RN(n1422), .Q(npc2[29]), .QN(
        net3429) );
  DFFR_X1 \npc2_reg[30]  ( .D(n232), .CK(Clk), .RN(n1422), .Q(npc2[30]), .QN(
        net3430) );
  DFFR_X1 \PC_reg[0]  ( .D(n231), .CK(Clk), .RN(n1418), .Q(PC[0]), .QN(net3464) );
  DFFR_X1 \PC_reg[1]  ( .D(n230), .CK(Clk), .RN(n1420), .Q(PC[1]), .QN(net3465) );
  DFFR_X1 \PC_reg[5]  ( .D(n226), .CK(Clk), .RN(n1419), .Q(PC[5]), .QN(net3469) );
  DFFR_X1 \PC_reg[6]  ( .D(n225), .CK(Clk), .RN(n1418), .Q(PC[6]), .QN(net3470) );
  DFFR_X1 \PC_reg[8]  ( .D(n223), .CK(Clk), .RN(n1418), .Q(PC[8]), .QN(net3472) );
  DFFR_X1 \PC_reg[10]  ( .D(n221), .CK(Clk), .RN(n1418), .Q(PC[10]), .QN(
        net3474) );
  DFFR_X1 \PC_reg[11]  ( .D(n220), .CK(Clk), .RN(n1419), .Q(PC[11]), .QN(
        net3475) );
  DFFR_X1 \PC_reg[12]  ( .D(n219), .CK(Clk), .RN(n1419), .Q(PC[12]), .QN(
        net3476) );
  DFFR_X1 \PC_reg[13]  ( .D(n218), .CK(Clk), .RN(n1419), .Q(PC[13]), .QN(
        net3477) );
  DFFR_X1 \PC_reg[14]  ( .D(n217), .CK(Clk), .RN(n1419), .Q(PC[14]), .QN(
        net3478) );
  DFFR_X1 \PC_reg[15]  ( .D(n216), .CK(Clk), .RN(n1419), .Q(PC[15]), .QN(
        net3479) );
  DFFR_X1 \PC_reg[16]  ( .D(n215), .CK(Clk), .RN(n1419), .Q(PC[16]), .QN(
        net3480) );
  DFFR_X1 \PC_reg[17]  ( .D(n214), .CK(Clk), .RN(n1423), .Q(PC[17]), .QN(
        net3481) );
  DFFR_X1 \PC_reg[18]  ( .D(n213), .CK(Clk), .RN(n1423), .Q(PC[18]), .QN(
        net3482) );
  DFFR_X1 \PC_reg[19]  ( .D(n212), .CK(Clk), .RN(n1423), .Q(PC[19]), .QN(
        net3483) );
  DFFR_X1 \PC_reg[20]  ( .D(n211), .CK(Clk), .RN(n1422), .Q(PC[20]), .QN(
        net3484) );
  DFFR_X1 \PC_reg[22]  ( .D(n209), .CK(Clk), .RN(n1422), .Q(PC[22]), .QN(
        net3486) );
  DFFR_X1 \PC_reg[23]  ( .D(n208), .CK(Clk), .RN(n1422), .Q(PC[23]), .QN(
        net3487) );
  DFFR_X1 \PC_reg[24]  ( .D(n207), .CK(Clk), .RN(n1418), .Q(PC[24]), .QN(
        net3488) );
  DFFR_X1 \PC_reg[25]  ( .D(n206), .CK(Clk), .RN(n1419), .Q(PC[25]), .QN(
        net3489) );
  DFFR_X1 \PC_reg[26]  ( .D(n205), .CK(Clk), .RN(n1419), .Q(PC[26]), .QN(
        net3490) );
  DFFR_X1 \PC_reg[27]  ( .D(n204), .CK(Clk), .RN(n1422), .Q(PC[27]), .QN(
        net3491) );
  DFFR_X1 \PC_reg[28]  ( .D(n203), .CK(Clk), .RN(n1422), .Q(PC[28]), .QN(
        net3492) );
  DFFR_X1 \PC_reg[29]  ( .D(n202), .CK(Clk), .RN(n1422), .Q(PC[29]), .QN(
        net3493) );
  DFFR_X1 \PC_reg[30]  ( .D(n201), .CK(Clk), .RN(n1422), .Q(PC[30]), .QN(
        net3494) );
  DFFR_X1 \IR_reg[7]  ( .D(n200), .CK(Clk), .RN(n1425), .Q(IR[7]), .QN(net3503) );
  DFFR_X1 \IR_reg[5]  ( .D(n199), .CK(Clk), .RN(n1425), .Q(IR[5]), .QN(net3501) );
  DFFR_X1 \IR_reg[3]  ( .D(n198), .CK(Clk), .RN(n1425), .Q(IR[3]), .QN(net3499) );
  DFFR_X1 \IR_reg[31]  ( .D(n197), .CK(Clk), .RN(n1425), .Q(IR[31]), .QN(
        net3527) );
  DFFR_X1 \IR_reg[29]  ( .D(n196), .CK(Clk), .RN(n1425), .Q(IR[29]), .QN(
        net3525) );
  DFFR_X1 \IR_reg[1]  ( .D(n195), .CK(Clk), .RN(n1425), .Q(IR[1]), .QN(net3497) );
  DFFR_X1 \IR_reg[26]  ( .D(n194), .CK(Clk), .RN(n1425), .Q(IR[26]), .QN(
        net3522) );
  DFFR_X1 \IR_reg[24]  ( .D(n193), .CK(Clk), .RN(n1425), .Q(IR[24]), .QN(
        net3520) );
  DFFR_X1 \IR_reg[22]  ( .D(n192), .CK(Clk), .RN(n1425), .Q(IR[22]), .QN(
        net3518) );
  DFFR_X1 \IR_reg[20]  ( .D(n191), .CK(Clk), .RN(n1425), .Q(IR[20]), .QN(
        net3516) );
  DFFR_X1 \IR_reg[18]  ( .D(n190), .CK(Clk), .RN(n1425), .Q(IR[18]), .QN(
        net3514) );
  DFFR_X1 \IR_reg[17]  ( .D(n189), .CK(Clk), .RN(n1424), .Q(IR[17]), .QN(
        net3513) );
  DFFR_X1 \IR_reg[15]  ( .D(n188), .CK(Clk), .RN(n1424), .Q(IR[15]), .QN(
        net3511) );
  DFFR_X1 \IR_reg[13]  ( .D(n187), .CK(Clk), .RN(n1424), .Q(IR[13]), .QN(
        net3509) );
  DFFR_X1 \IR_reg[11]  ( .D(n186), .CK(Clk), .RN(n1424), .Q(IR[11]), .QN(
        net3507) );
  DFFR_X1 \IR_reg[9]  ( .D(n185), .CK(Clk), .RN(n1424), .Q(IR[9]), .QN(net3505) );
  DFFR_X1 \IR_reg[8]  ( .D(n184), .CK(Clk), .RN(n1424), .Q(IR[8]), .QN(net3504) );
  DFFR_X1 \IR_reg[10]  ( .D(n183), .CK(Clk), .RN(n1424), .Q(IR[10]), .QN(
        net3506) );
  DFFR_X1 \IR_reg[12]  ( .D(n182), .CK(Clk), .RN(n1424), .Q(IR[12]), .QN(
        net3508) );
  DFFR_X1 \IR_reg[14]  ( .D(n181), .CK(Clk), .RN(n1424), .Q(IR[14]), .QN(
        net3510) );
  DFFR_X1 \IR_reg[16]  ( .D(n180), .CK(Clk), .RN(n1424), .Q(IR[16]), .QN(
        net3512) );
  DFFR_X1 \IR_reg[0]  ( .D(n179), .CK(Clk), .RN(n1424), .Q(IR[0]), .QN(net3496) );
  DFFR_X1 \IR_reg[19]  ( .D(n178), .CK(Clk), .RN(n1426), .Q(IR[19]), .QN(
        net3515) );
  DFFR_X1 \IR_reg[21]  ( .D(n177), .CK(Clk), .RN(n1426), .Q(IR[21]), .QN(
        net3517) );
  DFFR_X1 \IR_reg[23]  ( .D(n176), .CK(Clk), .RN(n1426), .Q(IR[23]), .QN(
        net3519) );
  DFFR_X1 \IR_reg[25]  ( .D(n175), .CK(Clk), .RN(n1426), .Q(IR[25]), .QN(
        net3521) );
  DFFR_X1 \IR_reg[27]  ( .D(n174), .CK(Clk), .RN(n1426), .Q(IR[27]), .QN(
        net3523) );
  DFFR_X1 \IR_reg[28]  ( .D(n173), .CK(Clk), .RN(n1426), .Q(IR[28]), .QN(
        net3524) );
  DFFR_X1 \IR_reg[30]  ( .D(n172), .CK(Clk), .RN(n1426), .Q(IR[30]), .QN(
        net3526) );
  DFFR_X1 \IR_reg[2]  ( .D(n171), .CK(Clk), .RN(n1426), .Q(IR[2]), .QN(net3498) );
  DFFR_X1 \IR_reg[4]  ( .D(n170), .CK(Clk), .RN(n1426), .Q(IR[4]), .QN(net3500) );
  DFFR_X1 \IR_reg[6]  ( .D(n169), .CK(Clk), .RN(n1426), .Q(IR[6]), .QN(net3502) );
  DFFR_X1 \PC_reg[4]  ( .D(n227), .CK(Clk), .RN(n1419), .Q(PC[4]), .QN(net3468) );
  DFFR_X1 \PC_reg[31]  ( .D(n295), .CK(Clk), .RN(n1422), .Q(PC[31]), .QN(
        net3495) );
  DFFR_X1 \PC_reg[9]  ( .D(n222), .CK(Clk), .RN(n1418), .Q(PC[9]), .QN(net3473) );
  DFFR_X1 \PC_reg[7]  ( .D(n224), .CK(Clk), .RN(n1418), .Q(PC[7]), .QN(net3471) );
  DFFR_X1 \PC_reg[3]  ( .D(n228), .CK(Clk), .RN(n1421), .Q(PC[3]), .QN(net3467) );
  DFFR_X1 \PC_reg[2]  ( .D(n229), .CK(Clk), .RN(n1421), .Q(PC[2]), .QN(net3466) );
  DFFR_X1 \PC_reg[21]  ( .D(n210), .CK(Clk), .RN(n1418), .Q(PC[21]), .QN(
        net3485) );
  datapath_reg_size32 DP_I ( .clk(Clk), .rst(n1418), .flush(n1225), .RF1(rd1_i), .RF2(rd2_i), .WF1(wr_i), .EN_regA(RegA_LATCH_EN_i), .EN_regB(RegB_LATCH_EN_i), .EN_regIMM(RegIMM_LATCH_EN_i), .EN_regALUOP(n1432), .EN_regRD1(en_RD1_i), 
        .EN_regNPC2(n1429), .S1(MUXA_SEL_i), .S2(MUXB_SEL_i), .EN_regRET(
        RETURN_REG_EN_i), .EN_regOUTALU(ALU_OUTREG_EN_i), .EN_regB2(B2_EN_i), 
        .EN_regRD2(en_RD2_i), .EN_regALU2(Alu_outreg2_en_i), .EN_regLMD(
        LMD_LATCH_EN_i), .EN_regRD3(en_RD3_i), .Sel_ret_alu(sel_alu_ret_i), 
        .Sel_alu_lmd(WB_MUX_SEL_i), .sel_31_rd(wb_mux_add_sel_i), .NPC(out_NPC), .IR_dp(IR), .comp_branch_i(comp_branch_dp), .immediate_branch(immediate), 
        .ADD_mem(dram_ADD), .DIN_mem(dram_DIN), .DOUT_mem(dram_DOUT) );
  mux21_N32_0 mux_pc ( .A(in_NPC), .B(pc_jump), .SEL(n1225), .Y(PC_BUS) );
  CU_HDW_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE21 CU_I ( 
        .Clk(Clk), .Rst(n1418), .IR_IN(iram_Dout), .flush(n1225), 
        .NPC1_LATCH_EN(NPC1_LATCH_EN_i), .NPC2_LATCH_EN(n1230), 
        .RegA_LATCH_EN(RegA_LATCH_EN_i), .RegB_LATCH_EN(RegB_LATCH_EN_i), 
        .RegAluOpCodeGen_EN(n1233), .RegIMM_LATCH_EN(RegIMM_LATCH_EN_i), 
        .Reg_RD1_EN(en_RD1_i), .RD1(rd1_i), .RD2(rd2_i), .B2_LATCH_EN(B2_EN_i), 
        .MUXA_SEL(MUXA_SEL_i), .MUXB_SEL(MUXB_SEL_i), .ALU_OUTREG_EN(
        ALU_OUTREG_EN_i), .RETURN_REG_EN(RETURN_REG_EN_i), .Reg_RD2_EN(
        en_RD2_i), .ALU_OUT2_SEL(sel_alu_ret_i), .LMD_LATCH_EN(LMD_LATCH_EN_i), 
        .Alu_outreg2_en(Alu_outreg2_en_i), .JUMP_en(JUMP_EN_i), .Reg_RD3_EN(
        en_RD3_i), .write_stop_if_branch(write_stop_if_branch_i), .WB_MUX_SEL(
        WB_MUX_SEL_i), .WB_MUX_ADD_SEL(wb_mux_add_sel_i), .WR(wr_cu) );
  DLX_IR_SIZE32_PC_SIZE32_DW01_add_0 add_351 ( .A(npc2), .B(immediate), .CI(
        1'b0), .SUM(pc_jump) );
  DLX_IR_SIZE32_PC_SIZE32_DW01_add_1 add_306 ( .A(PC), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0}), .CI(1'b0), .SUM(in_NPC) );
  DFFR_X1 \out_NPC_reg[31]  ( .D(n294), .CK(Clk), .RN(n1244), .Q(out_NPC[31]), 
        .QN(n1288) );
  DFFR_X1 \out_NPC_reg[30]  ( .D(n233), .CK(Clk), .RN(n1244), .Q(out_NPC[30]), 
        .QN(n1349) );
  DFFR_X1 \out_NPC_reg[29]  ( .D(n235), .CK(Clk), .RN(n1244), .Q(out_NPC[29]), 
        .QN(n1347) );
  DFFR_X1 \out_NPC_reg[28]  ( .D(n237), .CK(Clk), .RN(n1244), .Q(out_NPC[28]), 
        .QN(n1345) );
  DFFR_X1 \out_NPC_reg[27]  ( .D(n239), .CK(Clk), .RN(n1244), .Q(out_NPC[27]), 
        .QN(n1343) );
  DFFR_X1 \out_NPC_reg[26]  ( .D(n241), .CK(Clk), .RN(n1244), .Q(out_NPC[26]), 
        .QN(n1341) );
  DFFR_X1 \out_NPC_reg[25]  ( .D(n243), .CK(Clk), .RN(n1244), .Q(out_NPC[25]), 
        .QN(n1339) );
  DFFR_X1 \out_NPC_reg[24]  ( .D(n245), .CK(Clk), .RN(n1244), .Q(out_NPC[24]), 
        .QN(n1337) );
  DFFR_X1 \out_NPC_reg[23]  ( .D(n247), .CK(Clk), .RN(n1244), .Q(out_NPC[23]), 
        .QN(n1335) );
  DFFR_X1 \out_NPC_reg[22]  ( .D(n249), .CK(Clk), .RN(n1244), .Q(out_NPC[22]), 
        .QN(n1333) );
  DFFR_X1 \out_NPC_reg[21]  ( .D(n251), .CK(Clk), .RN(n1244), .Q(out_NPC[21]), 
        .QN(n1331) );
  DFFR_X1 \out_NPC_reg[20]  ( .D(n253), .CK(Clk), .RN(n1244), .Q(out_NPC[20]), 
        .QN(n1329) );
  DFFR_X1 \out_NPC_reg[19]  ( .D(n255), .CK(Clk), .RN(n1244), .Q(out_NPC[19]), 
        .QN(n1327) );
  DFFR_X1 \out_NPC_reg[18]  ( .D(n257), .CK(Clk), .RN(n1244), .Q(out_NPC[18]), 
        .QN(n1325) );
  DFFR_X1 \out_NPC_reg[17]  ( .D(n259), .CK(Clk), .RN(n1244), .Q(out_NPC[17]), 
        .QN(n1323) );
  DFFR_X1 \out_NPC_reg[16]  ( .D(n261), .CK(Clk), .RN(n1244), .Q(out_NPC[16]), 
        .QN(n1321) );
  DFFR_X1 \out_NPC_reg[15]  ( .D(n263), .CK(Clk), .RN(n1244), .Q(out_NPC[15]), 
        .QN(n1319) );
  DFFR_X1 \out_NPC_reg[14]  ( .D(n265), .CK(Clk), .RN(n1244), .Q(out_NPC[14]), 
        .QN(n1317) );
  DFFR_X1 \out_NPC_reg[13]  ( .D(n267), .CK(Clk), .RN(n1244), .Q(out_NPC[13]), 
        .QN(n1315) );
  DFFR_X1 \out_NPC_reg[12]  ( .D(n269), .CK(Clk), .RN(n1244), .Q(out_NPC[12]), 
        .QN(n1313) );
  DFFR_X1 \out_NPC_reg[11]  ( .D(n271), .CK(Clk), .RN(n1244), .Q(out_NPC[11]), 
        .QN(n1311) );
  DFFR_X1 \out_NPC_reg[10]  ( .D(n273), .CK(Clk), .RN(n1244), .Q(out_NPC[10]), 
        .QN(n1309) );
  DFFR_X1 \out_NPC_reg[9]  ( .D(n275), .CK(Clk), .RN(n1244), .Q(out_NPC[9]), 
        .QN(n1307) );
  DFFR_X1 \out_NPC_reg[8]  ( .D(n277), .CK(Clk), .RN(n1244), .Q(out_NPC[8]), 
        .QN(n1305) );
  DFFR_X1 \out_NPC_reg[7]  ( .D(n279), .CK(Clk), .RN(n1244), .Q(out_NPC[7]), 
        .QN(n1303) );
  DFFR_X1 \out_NPC_reg[6]  ( .D(n281), .CK(Clk), .RN(n1244), .Q(out_NPC[6]), 
        .QN(n1301) );
  DFFR_X1 \out_NPC_reg[5]  ( .D(n283), .CK(Clk), .RN(n1244), .Q(out_NPC[5]), 
        .QN(n1299) );
  DFFR_X1 \out_NPC_reg[4]  ( .D(n285), .CK(Clk), .RN(n1244), .Q(out_NPC[4]), 
        .QN(n1297) );
  DFFR_X1 \out_NPC_reg[3]  ( .D(n287), .CK(Clk), .RN(n1244), .Q(out_NPC[3]), 
        .QN(n1295) );
  DFFR_X1 \out_NPC_reg[2]  ( .D(n289), .CK(Clk), .RN(n1244), .Q(out_NPC[2]), 
        .QN(n1293) );
  DFFR_X1 \out_NPC_reg[1]  ( .D(n291), .CK(Clk), .RN(n1244), .Q(out_NPC[1]), 
        .QN(n1291) );
  DFFR_X1 \out_NPC_reg[0]  ( .D(n292), .CK(Clk), .RN(n1244), .Q(out_NPC[0]), 
        .QN(n1286) );
  OR2_X1 U1863 ( .A1(net3485), .A2(n1417), .ZN(n1415) );
  NAND2_X1 U1864 ( .A1(n1415), .A2(n1372), .ZN(n210) );
  OR2_X2 U1865 ( .A1(JUMP_EN_i), .A2(comp_branch_dp), .ZN(n1225) );
  BUF_X4 U1866 ( .A(NPC1_LATCH_EN_i), .Z(n1417) );
  BUF_X4 U1867 ( .A(NPC1_LATCH_EN_i), .Z(n1416) );
  INV_X1 U1868 ( .A(n1432), .ZN(n1430) );
  INV_X1 U1869 ( .A(n1435), .ZN(n1431) );
  BUF_X1 U1870 ( .A(n1427), .Z(n1432) );
  BUF_X1 U1871 ( .A(n1427), .Z(n1433) );
  BUF_X1 U1872 ( .A(n1428), .Z(n1434) );
  BUF_X1 U1873 ( .A(n1428), .Z(n1435) );
  BUF_X1 U1874 ( .A(n1230), .Z(n1429) );
  BUF_X1 U1875 ( .A(n1233), .Z(n1427) );
  BUF_X1 U1876 ( .A(n1233), .Z(n1428) );
  BUF_X1 U1877 ( .A(n1238), .Z(n1424) );
  BUF_X1 U1878 ( .A(n1238), .Z(n1425) );
  BUF_X1 U1879 ( .A(n1238), .Z(n1426) );
  OAI21_X1 U1880 ( .B1(n1416), .B2(n1349), .A(n1350), .ZN(n233) );
  NAND2_X1 U1881 ( .A1(in_NPC[30]), .A2(n1416), .ZN(n1350) );
  OAI21_X1 U1882 ( .B1(n1416), .B2(n1297), .A(n1298), .ZN(n285) );
  NAND2_X1 U1883 ( .A1(in_NPC[4]), .A2(n1416), .ZN(n1298) );
  OAI21_X1 U1884 ( .B1(n1416), .B2(n1317), .A(n1318), .ZN(n265) );
  NAND2_X1 U1885 ( .A1(in_NPC[14]), .A2(n1416), .ZN(n1318) );
  OAI21_X1 U1886 ( .B1(n1416), .B2(n1321), .A(n1322), .ZN(n261) );
  NAND2_X1 U1887 ( .A1(in_NPC[16]), .A2(n1416), .ZN(n1322) );
  OAI21_X1 U1888 ( .B1(n1416), .B2(n1337), .A(n1338), .ZN(n245) );
  NAND2_X1 U1889 ( .A1(in_NPC[24]), .A2(n1416), .ZN(n1338) );
  OAI21_X1 U1890 ( .B1(n1417), .B2(n1299), .A(n1300), .ZN(n283) );
  NAND2_X1 U1891 ( .A1(in_NPC[5]), .A2(n1416), .ZN(n1300) );
  OAI21_X1 U1892 ( .B1(n1417), .B2(n1307), .A(n1308), .ZN(n275) );
  NAND2_X1 U1893 ( .A1(in_NPC[9]), .A2(n1416), .ZN(n1308) );
  OAI21_X1 U1894 ( .B1(n1417), .B2(n1327), .A(n1328), .ZN(n255) );
  NAND2_X1 U1895 ( .A1(in_NPC[19]), .A2(n1416), .ZN(n1328) );
  OAI21_X1 U1896 ( .B1(n1417), .B2(n1335), .A(n1336), .ZN(n247) );
  NAND2_X1 U1897 ( .A1(in_NPC[23]), .A2(n1416), .ZN(n1336) );
  OAI21_X1 U1898 ( .B1(n1417), .B2(n1339), .A(n1340), .ZN(n243) );
  NAND2_X1 U1899 ( .A1(in_NPC[25]), .A2(n1416), .ZN(n1340) );
  OAI21_X1 U1900 ( .B1(n1417), .B2(n1347), .A(n1348), .ZN(n235) );
  NAND2_X1 U1901 ( .A1(in_NPC[29]), .A2(n1416), .ZN(n1348) );
  OAI21_X1 U1902 ( .B1(n1416), .B2(n1301), .A(n1302), .ZN(n281) );
  NAND2_X1 U1903 ( .A1(in_NPC[6]), .A2(n1417), .ZN(n1302) );
  OAI21_X1 U1904 ( .B1(n1416), .B2(n1305), .A(n1306), .ZN(n277) );
  NAND2_X1 U1905 ( .A1(in_NPC[8]), .A2(n1417), .ZN(n1306) );
  OAI21_X1 U1906 ( .B1(n1416), .B2(n1309), .A(n1310), .ZN(n273) );
  NAND2_X1 U1907 ( .A1(in_NPC[10]), .A2(n1417), .ZN(n1310) );
  OAI21_X1 U1908 ( .B1(n1416), .B2(n1313), .A(n1314), .ZN(n269) );
  NAND2_X1 U1909 ( .A1(in_NPC[12]), .A2(n1417), .ZN(n1314) );
  OAI21_X1 U1910 ( .B1(n1416), .B2(n1325), .A(n1326), .ZN(n257) );
  NAND2_X1 U1911 ( .A1(in_NPC[18]), .A2(n1417), .ZN(n1326) );
  OAI21_X1 U1912 ( .B1(n1416), .B2(n1329), .A(n1330), .ZN(n253) );
  NAND2_X1 U1913 ( .A1(in_NPC[20]), .A2(n1417), .ZN(n1330) );
  OAI21_X1 U1914 ( .B1(n1416), .B2(n1333), .A(n1334), .ZN(n249) );
  NAND2_X1 U1915 ( .A1(in_NPC[22]), .A2(n1417), .ZN(n1334) );
  OAI21_X1 U1916 ( .B1(n1416), .B2(n1341), .A(n1342), .ZN(n241) );
  NAND2_X1 U1917 ( .A1(in_NPC[26]), .A2(n1417), .ZN(n1342) );
  OAI21_X1 U1918 ( .B1(n1416), .B2(n1345), .A(n1346), .ZN(n237) );
  NAND2_X1 U1919 ( .A1(in_NPC[28]), .A2(n1417), .ZN(n1346) );
  OAI21_X1 U1920 ( .B1(n1416), .B2(n1288), .A(n1289), .ZN(n294) );
  NAND2_X1 U1921 ( .A1(in_NPC[31]), .A2(n1417), .ZN(n1289) );
  OAI21_X1 U1922 ( .B1(n1417), .B2(n1293), .A(n1294), .ZN(n289) );
  NAND2_X1 U1923 ( .A1(in_NPC[2]), .A2(n1417), .ZN(n1294) );
  OAI21_X1 U1924 ( .B1(n1417), .B2(n1295), .A(n1296), .ZN(n287) );
  NAND2_X1 U1925 ( .A1(in_NPC[3]), .A2(n1417), .ZN(n1296) );
  OAI21_X1 U1926 ( .B1(n1417), .B2(n1303), .A(n1304), .ZN(n279) );
  NAND2_X1 U1927 ( .A1(in_NPC[7]), .A2(n1417), .ZN(n1304) );
  OAI21_X1 U1928 ( .B1(n1417), .B2(n1311), .A(n1312), .ZN(n271) );
  NAND2_X1 U1929 ( .A1(in_NPC[11]), .A2(n1417), .ZN(n1312) );
  OAI21_X1 U1930 ( .B1(n1417), .B2(n1315), .A(n1316), .ZN(n267) );
  NAND2_X1 U1931 ( .A1(in_NPC[13]), .A2(n1417), .ZN(n1316) );
  OAI21_X1 U1932 ( .B1(n1417), .B2(n1319), .A(n1320), .ZN(n263) );
  NAND2_X1 U1933 ( .A1(in_NPC[15]), .A2(n1417), .ZN(n1320) );
  OAI21_X1 U1934 ( .B1(n1417), .B2(n1323), .A(n1324), .ZN(n259) );
  NAND2_X1 U1935 ( .A1(in_NPC[17]), .A2(n1417), .ZN(n1324) );
  OAI21_X1 U1936 ( .B1(n1417), .B2(n1331), .A(n1332), .ZN(n251) );
  NAND2_X1 U1937 ( .A1(in_NPC[21]), .A2(n1417), .ZN(n1332) );
  OAI21_X1 U1938 ( .B1(n1417), .B2(n1343), .A(n1344), .ZN(n239) );
  NAND2_X1 U1939 ( .A1(in_NPC[27]), .A2(n1417), .ZN(n1344) );
  AND2_X1 U1940 ( .A1(n1423), .A2(n1414), .ZN(n1238) );
  NOR2_X1 U1941 ( .A1(JUMP_EN_i), .A2(comp_branch_dp), .ZN(n1414) );
  NAND2_X1 U1942 ( .A1(PC_BUS[21]), .A2(n1416), .ZN(n1372) );
  OAI21_X1 U1943 ( .B1(net3494), .B2(n1416), .A(n1381), .ZN(n201) );
  NAND2_X1 U1944 ( .A1(PC_BUS[30]), .A2(n1416), .ZN(n1381) );
  OAI21_X1 U1945 ( .B1(net3493), .B2(n1416), .A(n1380), .ZN(n202) );
  NAND2_X1 U1946 ( .A1(PC_BUS[29]), .A2(n1416), .ZN(n1380) );
  OAI21_X1 U1947 ( .B1(net3492), .B2(n1416), .A(n1379), .ZN(n203) );
  NAND2_X1 U1948 ( .A1(PC_BUS[28]), .A2(n1417), .ZN(n1379) );
  OAI21_X1 U1949 ( .B1(net3491), .B2(n1416), .A(n1378), .ZN(n204) );
  NAND2_X1 U1950 ( .A1(PC_BUS[27]), .A2(n1417), .ZN(n1378) );
  OAI21_X1 U1951 ( .B1(net3490), .B2(n1416), .A(n1377), .ZN(n205) );
  NAND2_X1 U1952 ( .A1(PC_BUS[26]), .A2(n1416), .ZN(n1377) );
  OAI21_X1 U1953 ( .B1(net3489), .B2(n1417), .A(n1376), .ZN(n206) );
  NAND2_X1 U1954 ( .A1(PC_BUS[25]), .A2(n1417), .ZN(n1376) );
  OAI21_X1 U1955 ( .B1(net3488), .B2(n1417), .A(n1375), .ZN(n207) );
  NAND2_X1 U1956 ( .A1(PC_BUS[24]), .A2(n1416), .ZN(n1375) );
  OAI21_X1 U1957 ( .B1(net3487), .B2(n1417), .A(n1374), .ZN(n208) );
  NAND2_X1 U1958 ( .A1(PC_BUS[23]), .A2(n1416), .ZN(n1374) );
  OAI21_X1 U1959 ( .B1(net3486), .B2(n1417), .A(n1373), .ZN(n209) );
  NAND2_X1 U1960 ( .A1(PC_BUS[22]), .A2(n1416), .ZN(n1373) );
  OAI21_X1 U1961 ( .B1(net3484), .B2(n1417), .A(n1371), .ZN(n211) );
  NAND2_X1 U1962 ( .A1(PC_BUS[20]), .A2(n1416), .ZN(n1371) );
  OAI21_X1 U1963 ( .B1(net3483), .B2(n1417), .A(n1370), .ZN(n212) );
  NAND2_X1 U1964 ( .A1(PC_BUS[19]), .A2(n1416), .ZN(n1370) );
  OAI21_X1 U1965 ( .B1(net3482), .B2(n1417), .A(n1369), .ZN(n213) );
  NAND2_X1 U1966 ( .A1(PC_BUS[18]), .A2(n1416), .ZN(n1369) );
  OAI21_X1 U1967 ( .B1(net3481), .B2(n1416), .A(n1368), .ZN(n214) );
  NAND2_X1 U1968 ( .A1(PC_BUS[17]), .A2(n1416), .ZN(n1368) );
  OAI21_X1 U1969 ( .B1(net3480), .B2(n1416), .A(n1367), .ZN(n215) );
  NAND2_X1 U1970 ( .A1(PC_BUS[16]), .A2(n1416), .ZN(n1367) );
  OAI21_X1 U1971 ( .B1(net3479), .B2(n1417), .A(n1366), .ZN(n216) );
  NAND2_X1 U1972 ( .A1(PC_BUS[15]), .A2(n1416), .ZN(n1366) );
  OAI21_X1 U1973 ( .B1(net3478), .B2(n1417), .A(n1365), .ZN(n217) );
  NAND2_X1 U1974 ( .A1(PC_BUS[14]), .A2(n1417), .ZN(n1365) );
  OAI21_X1 U1975 ( .B1(net3477), .B2(n1417), .A(n1364), .ZN(n218) );
  NAND2_X1 U1976 ( .A1(PC_BUS[13]), .A2(n1417), .ZN(n1364) );
  OAI21_X1 U1977 ( .B1(net3476), .B2(n1416), .A(n1363), .ZN(n219) );
  NAND2_X1 U1978 ( .A1(PC_BUS[12]), .A2(n1417), .ZN(n1363) );
  OAI21_X1 U1979 ( .B1(net3475), .B2(n1417), .A(n1362), .ZN(n220) );
  NAND2_X1 U1980 ( .A1(PC_BUS[11]), .A2(n1417), .ZN(n1362) );
  OAI21_X1 U1981 ( .B1(net3474), .B2(n1416), .A(n1361), .ZN(n221) );
  NAND2_X1 U1982 ( .A1(PC_BUS[10]), .A2(n1416), .ZN(n1361) );
  OAI21_X1 U1983 ( .B1(net3464), .B2(n1416), .A(n1351), .ZN(n231) );
  NAND2_X1 U1984 ( .A1(PC_BUS[0]), .A2(n1417), .ZN(n1351) );
  OAI21_X1 U1985 ( .B1(net3466), .B2(n1417), .A(n1353), .ZN(n229) );
  NAND2_X1 U1986 ( .A1(PC_BUS[2]), .A2(n1417), .ZN(n1353) );
  OAI21_X1 U1987 ( .B1(net3465), .B2(n1417), .A(n1352), .ZN(n230) );
  NAND2_X1 U1988 ( .A1(PC_BUS[1]), .A2(n1417), .ZN(n1352) );
  OAI21_X1 U1989 ( .B1(net3467), .B2(n1416), .A(n1354), .ZN(n228) );
  NAND2_X1 U1990 ( .A1(PC_BUS[3]), .A2(n1416), .ZN(n1354) );
  OAI21_X1 U1991 ( .B1(net3471), .B2(n1417), .A(n1358), .ZN(n224) );
  NAND2_X1 U1992 ( .A1(PC_BUS[7]), .A2(n1416), .ZN(n1358) );
  OAI21_X1 U1993 ( .B1(net3473), .B2(n1416), .A(n1360), .ZN(n222) );
  NAND2_X1 U1994 ( .A1(PC_BUS[9]), .A2(n1416), .ZN(n1360) );
  OAI21_X1 U1995 ( .B1(net3468), .B2(n1417), .A(n1355), .ZN(n227) );
  NAND2_X1 U1996 ( .A1(PC_BUS[4]), .A2(n1417), .ZN(n1355) );
  OAI21_X1 U1997 ( .B1(net3472), .B2(n1417), .A(n1359), .ZN(n223) );
  NAND2_X1 U1998 ( .A1(PC_BUS[8]), .A2(n1416), .ZN(n1359) );
  OAI21_X1 U1999 ( .B1(net3470), .B2(n1416), .A(n1357), .ZN(n225) );
  NAND2_X1 U2000 ( .A1(PC_BUS[6]), .A2(n1416), .ZN(n1357) );
  OAI21_X1 U2001 ( .B1(net3469), .B2(n1416), .A(n1356), .ZN(n226) );
  NAND2_X1 U2002 ( .A1(PC_BUS[5]), .A2(n1417), .ZN(n1356) );
  OAI21_X1 U2003 ( .B1(net3495), .B2(n1416), .A(n1287), .ZN(n295) );
  NAND2_X1 U2004 ( .A1(PC_BUS[31]), .A2(n1417), .ZN(n1287) );
  OAI22_X1 U2005 ( .A1(n1431), .A2(n1325), .B1(n1429), .B2(net3418), .ZN(n256)
         );
  OAI22_X1 U2006 ( .A1(n1431), .A2(n1323), .B1(n1429), .B2(net3417), .ZN(n258)
         );
  OAI22_X1 U2007 ( .A1(n1431), .A2(n1321), .B1(n1429), .B2(net3416), .ZN(n260)
         );
  OAI22_X1 U2008 ( .A1(n1431), .A2(n1319), .B1(n1429), .B2(net3415), .ZN(n262)
         );
  OAI22_X1 U2009 ( .A1(n1431), .A2(n1317), .B1(n1429), .B2(net3414), .ZN(n264)
         );
  OAI22_X1 U2010 ( .A1(n1431), .A2(n1315), .B1(n1429), .B2(net3413), .ZN(n266)
         );
  OAI22_X1 U2011 ( .A1(n1431), .A2(n1313), .B1(n1429), .B2(net3412), .ZN(n268)
         );
  OAI22_X1 U2012 ( .A1(n1431), .A2(n1311), .B1(n1429), .B2(net3411), .ZN(n270)
         );
  OAI22_X1 U2013 ( .A1(n1431), .A2(n1307), .B1(n1429), .B2(net3409), .ZN(n274)
         );
  OAI22_X1 U2014 ( .A1(n1431), .A2(n1305), .B1(n1429), .B2(net3408), .ZN(n276)
         );
  OAI22_X1 U2015 ( .A1(n1431), .A2(n1303), .B1(n1429), .B2(net3407), .ZN(n278)
         );
  OAI22_X1 U2016 ( .A1(n1431), .A2(n1301), .B1(n1429), .B2(net3406), .ZN(n280)
         );
  OAI22_X1 U2017 ( .A1(n1431), .A2(n1299), .B1(n1429), .B2(net3405), .ZN(n282)
         );
  OAI22_X1 U2018 ( .A1(n1431), .A2(n1297), .B1(n1429), .B2(net3404), .ZN(n284)
         );
  OAI22_X1 U2019 ( .A1(n1431), .A2(n1295), .B1(n1429), .B2(net3403), .ZN(n286)
         );
  OAI22_X1 U2020 ( .A1(n1431), .A2(n1293), .B1(n1429), .B2(net3402), .ZN(n288)
         );
  OAI22_X1 U2021 ( .A1(n1431), .A2(n1291), .B1(n1429), .B2(net3401), .ZN(n290)
         );
  OAI22_X1 U2022 ( .A1(n1431), .A2(n1288), .B1(n1429), .B2(net3431), .ZN(n293)
         );
  OAI22_X1 U2023 ( .A1(n1431), .A2(n1286), .B1(n1429), .B2(net3400), .ZN(n296)
         );
  OAI22_X1 U2024 ( .A1(n1430), .A2(n1331), .B1(n1432), .B2(net3421), .ZN(n250)
         );
  OAI22_X1 U2025 ( .A1(n1430), .A2(n1329), .B1(n1432), .B2(net3420), .ZN(n252)
         );
  OAI22_X1 U2026 ( .A1(n1431), .A2(n1327), .B1(n1432), .B2(net3419), .ZN(n254)
         );
  OAI22_X1 U2027 ( .A1(n1430), .A2(n1349), .B1(n1434), .B2(net3430), .ZN(n232)
         );
  OAI22_X1 U2028 ( .A1(n1430), .A2(n1347), .B1(n1434), .B2(net3429), .ZN(n234)
         );
  OAI22_X1 U2029 ( .A1(n1430), .A2(n1345), .B1(n1434), .B2(net3428), .ZN(n236)
         );
  OAI22_X1 U2030 ( .A1(n1430), .A2(n1343), .B1(n1434), .B2(net3427), .ZN(n238)
         );
  OAI22_X1 U2031 ( .A1(n1430), .A2(n1341), .B1(n1433), .B2(net3426), .ZN(n240)
         );
  OAI22_X1 U2032 ( .A1(n1430), .A2(n1339), .B1(n1433), .B2(net3425), .ZN(n242)
         );
  OAI22_X1 U2033 ( .A1(n1430), .A2(n1337), .B1(n1433), .B2(net3424), .ZN(n244)
         );
  OAI22_X1 U2034 ( .A1(n1430), .A2(n1335), .B1(n1433), .B2(net3423), .ZN(n246)
         );
  OAI22_X1 U2035 ( .A1(n1430), .A2(n1333), .B1(n1433), .B2(net3422), .ZN(n248)
         );
  OAI22_X1 U2036 ( .A1(n1431), .A2(n1309), .B1(n1434), .B2(net3410), .ZN(n272)
         );
  OAI21_X1 U2037 ( .B1(n1416), .B2(n1291), .A(n1292), .ZN(n291) );
  NAND2_X1 U2038 ( .A1(in_NPC[1]), .A2(n1416), .ZN(n1292) );
  OAI21_X1 U2039 ( .B1(n1417), .B2(n1286), .A(n1290), .ZN(n292) );
  NAND2_X1 U2040 ( .A1(in_NPC[0]), .A2(n1417), .ZN(n1290) );
  OAI21_X1 U2041 ( .B1(net3502), .B2(n1417), .A(n1413), .ZN(n169) );
  NAND2_X1 U2042 ( .A1(iram_Dout[6]), .A2(n1417), .ZN(n1413) );
  OAI21_X1 U2043 ( .B1(net3500), .B2(n1417), .A(n1412), .ZN(n170) );
  NAND2_X1 U2044 ( .A1(iram_Dout[4]), .A2(n1416), .ZN(n1412) );
  OAI21_X1 U2045 ( .B1(net3498), .B2(n1417), .A(n1411), .ZN(n171) );
  NAND2_X1 U2046 ( .A1(iram_Dout[2]), .A2(n1417), .ZN(n1411) );
  OAI21_X1 U2047 ( .B1(net3526), .B2(n1417), .A(n1410), .ZN(n172) );
  NAND2_X1 U2048 ( .A1(iram_Dout[30]), .A2(n1416), .ZN(n1410) );
  OAI21_X1 U2049 ( .B1(net3524), .B2(n1416), .A(n1409), .ZN(n173) );
  NAND2_X1 U2050 ( .A1(iram_Dout[28]), .A2(n1416), .ZN(n1409) );
  OAI21_X1 U2051 ( .B1(net3523), .B2(n1416), .A(n1408), .ZN(n174) );
  NAND2_X1 U2052 ( .A1(iram_Dout[27]), .A2(n1416), .ZN(n1408) );
  OAI21_X1 U2053 ( .B1(net3521), .B2(n1416), .A(n1407), .ZN(n175) );
  NAND2_X1 U2054 ( .A1(iram_Dout[25]), .A2(n1416), .ZN(n1407) );
  OAI21_X1 U2055 ( .B1(net3519), .B2(n1416), .A(n1406), .ZN(n176) );
  NAND2_X1 U2056 ( .A1(iram_Dout[23]), .A2(n1416), .ZN(n1406) );
  OAI21_X1 U2057 ( .B1(net3517), .B2(n1417), .A(n1405), .ZN(n177) );
  NAND2_X1 U2058 ( .A1(iram_Dout[21]), .A2(n1417), .ZN(n1405) );
  OAI21_X1 U2059 ( .B1(net3515), .B2(n1416), .A(n1404), .ZN(n178) );
  NAND2_X1 U2060 ( .A1(iram_Dout[19]), .A2(n1416), .ZN(n1404) );
  OAI21_X1 U2061 ( .B1(net3496), .B2(n1416), .A(n1403), .ZN(n179) );
  NAND2_X1 U2062 ( .A1(iram_Dout[0]), .A2(n1416), .ZN(n1403) );
  OAI21_X1 U2063 ( .B1(net3512), .B2(n1417), .A(n1402), .ZN(n180) );
  NAND2_X1 U2064 ( .A1(iram_Dout[16]), .A2(n1416), .ZN(n1402) );
  OAI21_X1 U2065 ( .B1(net3510), .B2(n1417), .A(n1401), .ZN(n181) );
  NAND2_X1 U2066 ( .A1(iram_Dout[14]), .A2(n1417), .ZN(n1401) );
  OAI21_X1 U2067 ( .B1(net3508), .B2(n1417), .A(n1400), .ZN(n182) );
  NAND2_X1 U2068 ( .A1(iram_Dout[12]), .A2(n1417), .ZN(n1400) );
  OAI21_X1 U2069 ( .B1(net3506), .B2(n1416), .A(n1399), .ZN(n183) );
  NAND2_X1 U2070 ( .A1(iram_Dout[10]), .A2(n1417), .ZN(n1399) );
  OAI21_X1 U2071 ( .B1(net3504), .B2(n1416), .A(n1398), .ZN(n184) );
  NAND2_X1 U2072 ( .A1(iram_Dout[8]), .A2(n1416), .ZN(n1398) );
  OAI21_X1 U2073 ( .B1(net3505), .B2(n1417), .A(n1397), .ZN(n185) );
  NAND2_X1 U2074 ( .A1(iram_Dout[9]), .A2(n1417), .ZN(n1397) );
  OAI21_X1 U2075 ( .B1(net3507), .B2(n1417), .A(n1396), .ZN(n186) );
  NAND2_X1 U2076 ( .A1(iram_Dout[11]), .A2(n1416), .ZN(n1396) );
  OAI21_X1 U2077 ( .B1(net3509), .B2(n1416), .A(n1395), .ZN(n187) );
  NAND2_X1 U2078 ( .A1(iram_Dout[13]), .A2(n1416), .ZN(n1395) );
  OAI21_X1 U2079 ( .B1(net3511), .B2(n1416), .A(n1394), .ZN(n188) );
  NAND2_X1 U2080 ( .A1(iram_Dout[15]), .A2(n1416), .ZN(n1394) );
  OAI21_X1 U2081 ( .B1(net3513), .B2(n1416), .A(n1393), .ZN(n189) );
  NAND2_X1 U2082 ( .A1(iram_Dout[17]), .A2(n1417), .ZN(n1393) );
  OAI21_X1 U2083 ( .B1(net3514), .B2(n1416), .A(n1392), .ZN(n190) );
  NAND2_X1 U2084 ( .A1(iram_Dout[18]), .A2(n1417), .ZN(n1392) );
  OAI21_X1 U2085 ( .B1(net3516), .B2(n1417), .A(n1391), .ZN(n191) );
  NAND2_X1 U2086 ( .A1(iram_Dout[20]), .A2(n1417), .ZN(n1391) );
  OAI21_X1 U2087 ( .B1(net3518), .B2(n1416), .A(n1390), .ZN(n192) );
  NAND2_X1 U2088 ( .A1(iram_Dout[22]), .A2(n1417), .ZN(n1390) );
  OAI21_X1 U2089 ( .B1(net3520), .B2(n1416), .A(n1389), .ZN(n193) );
  NAND2_X1 U2090 ( .A1(iram_Dout[24]), .A2(n1417), .ZN(n1389) );
  OAI21_X1 U2091 ( .B1(net3522), .B2(n1416), .A(n1388), .ZN(n194) );
  NAND2_X1 U2092 ( .A1(iram_Dout[26]), .A2(n1416), .ZN(n1388) );
  OAI21_X1 U2093 ( .B1(net3497), .B2(n1417), .A(n1387), .ZN(n195) );
  NAND2_X1 U2094 ( .A1(iram_Dout[1]), .A2(n1417), .ZN(n1387) );
  OAI21_X1 U2095 ( .B1(net3525), .B2(n1416), .A(n1386), .ZN(n196) );
  NAND2_X1 U2096 ( .A1(iram_Dout[29]), .A2(n1417), .ZN(n1386) );
  OAI21_X1 U2097 ( .B1(net3527), .B2(n1417), .A(n1385), .ZN(n197) );
  NAND2_X1 U2098 ( .A1(iram_Dout[31]), .A2(n1416), .ZN(n1385) );
  OAI21_X1 U2099 ( .B1(net3499), .B2(n1417), .A(n1384), .ZN(n198) );
  NAND2_X1 U2100 ( .A1(iram_Dout[3]), .A2(n1417), .ZN(n1384) );
  OAI21_X1 U2101 ( .B1(net3501), .B2(n1416), .A(n1383), .ZN(n199) );
  NAND2_X1 U2102 ( .A1(iram_Dout[5]), .A2(n1416), .ZN(n1383) );
  OAI21_X1 U2103 ( .B1(net3503), .B2(n1417), .A(n1382), .ZN(n200) );
  NAND2_X1 U2104 ( .A1(iram_Dout[7]), .A2(n1416), .ZN(n1382) );
  BUF_X1 U2105 ( .A(n1244), .Z(n1418) );
  NOR2_X1 U2106 ( .A1(write_stop_if_branch_i), .A2(n1284), .ZN(wr_i) );
  INV_X1 U2107 ( .A(wr_cu), .ZN(n1284) );
  CLKBUF_X1 U2108 ( .A(n1244), .Z(n1419) );
  CLKBUF_X1 U2109 ( .A(n1244), .Z(n1420) );
  CLKBUF_X1 U2110 ( .A(n1244), .Z(n1421) );
  CLKBUF_X1 U2111 ( .A(n1244), .Z(n1422) );
  CLKBUF_X1 U2112 ( .A(n1244), .Z(n1423) );
endmodule

