LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.numeric_std.all;
USE IEEE.std_logic_unsigned.all;
ENTITY DUT_handler IS
PORT(
  CLOCK_50:BUFFER STD_LOGIC;
OUTPUT_VALID,RD_ACK,WR_ACK,MEM_WRITTEN,MEM_READ,START_ACK :IN STD_LOGIC;
RESET, RD_REQ,WR_REQ,READ_READY,ENABLE_GENERATORE,START: BUFFER STD_LOGIC
);  
END ENTITY DUT_handler;
ARCHITECTURE BEH OF DUT_handler IS
  
  CONSTANT PERIODO : TIME := 20 ns;
  CONSTANT RESET_TIME : TIME := 45 ns;

  COMPONENT COUNTER_NBIT IS
GENERIC (N:INTEGER);
PORT(
EN_COUNT, LOAD_COUNT,CLK,RESET	: IN STD_LOGIC;	--abilita conta, carica dato da cui iniziare a contare
COUNT_IN	:	IN STD_LOGIC_VECTOR((N-1) DOWNTO 0);	--dato da caricare in parallelo
COUNT_OUT	:	OUT STD_LOGIC_VECTOR((N-1) DOWNTO 0);
TC	:	OUT STD_LOGIC	--terminal count
);
END COMPONENT;

 SIGNAL TOTALE_SCRITTURE:INTEGER;
 SIGNAL WRITE_FLAG,READ_FLAG:STD_LOGIC;
  BEGIN
 
GENERA_WRITE: PROCESS(CLOCK_50,RESET,WR_ACK,WRITE_FLAG)
VARIABLE FLAG_CONTA,TOT_CONTEGGI:INTEGER;
BEGIN

IF (RESET='0') THEN
  TOT_CONTEGGI:=0; FLAG_CONTA:=0; WR_REQ<='0'; ENABLE_GENERATORE<='0';TOTALE_SCRITTURE<=0;
ELSE

  IF (CLOCK_50'EVENT AND CLOCK_50='1') THEN
    IF(WRITE_FLAG='0') THEN
   IF (WR_ACK='1') THEN
WR_REQ<='0' ; ELSE  
IF (TOT_CONTEGGI<2**18+100) THEN 
FLAG_CONTA:=FLAG_CONTA+1;  
IF (FLAG_CONTA=5) THEN
IF(WR_ACK='0') THEN
TOT_CONTEGGI:=TOT_CONTEGGI+1; FLAG_CONTA:=0;WR_REQ<='1'; ENABLE_GENERATORE<='1'; 
TOTALE_SCRITTURE<=TOTALE_SCRITTURE+1;
ELSE
FLAG_CONTA:=FLAG_CONTA-1; 
END IF;  END IF;  END IF;  END IF;  END IF; END IF; END IF;
END PROCESS;


GENERA_START: PROCESS (CLOCK_50,RESET,TOTALE_SCRITTURE,START_ACK,START,READ_FLAG)
 VARIABLE FLAG:STD_LOGIC;
BEGIN
IF (RESET='0') THEN
    START<='0'; FLAG:='0';
ELSE
 IF (CLOCK_50'EVENT AND CLOCK_50='1') THEN 
  IF (READ_FLAG='0') THEN
  IF (START='0') THEN
  IF (START_ACK='0') THEN
  IF(TOTALE_SCRITTURE>2**17)THEN --ASPETTO 2^17 SCRITTURE PRIMA DI CHIEDERE LA LETTURA DELLA MEMORIA
  IF FLAG='0' THEN
  START<='1';
  FLAG:='1';
  END IF;
  END IF; 
  END IF;
ELSIF (START='1') THEN 
IF (START_ACK='1') THEN
START<='0';
     END IF;  END IF; END IF; END IF; END IF;
   END PROCESS;
   
GENERA_READ: PROCESS (CLOCK_50,RESET,RD_ACK,READ_FLAG,RD_REQ,MEM_WRITTEN)
BEGIN
IF (RESET='0') THEN
    RD_REQ<='0'; 
ELSE
 IF (CLOCK_50'EVENT AND CLOCK_50='1') THEN 
IF RD_REQ='0' THEN 
IF MEM_WRITTEN='1' THEN
  RD_REQ<='1';
ELSE RD_REQ<='0';
END IF;
ELSE 
IF RD_ACK='1' THEN
RD_REQ<='0'; 
ELSE RD_REQ<='1';
END IF; END IF; END IF; END IF; 
END PROCESS;
   
   
GESTORE_LETTURE: PROCESS(CLOCK_50,RESET,OUTPUT_VALID,READ_FLAG)
BEGIN  
IF (RESET='0') THEN
  READ_READY<='0';
  ELSE
 
    IF (CLOCK_50'EVENT AND CLOCK_50='1') THEN
  IF (READ_FLAG='0') THEN
  IF (OUTPUT_VALID='1') THEN
   READ_READY<='1';
ELSE READ_READY<='0';
   END  IF; END IF; END IF; END IF;
END PROCESS;   
   
GESTORE_PROCESSI_DUT_HANDLER:PROCESS(CLOCK_50,RESET,MEM_WRITTEN,MEM_READ)
BEGIN
IF (RESET='0') THEN
WRITE_FLAG<='0'; READ_FLAG<='0';
ELSIF(CLOCK_50'EVENT AND CLOCK_50='1') THEN
IF(MEM_WRITTEN='1') THEN WRITE_FLAG<='1';
END IF;
IF(MEM_READ='1') THEN READ_FLAG<='1';
END IF;  END IF;
END PROCESS;
   
   
RESET <= '0', '1' AFTER RESET_TIME;    
GENERATORE_CLOCK :PROCESS
   BEGIN
        CLOCK_50 <= '0';
        WAIT FOR PERIODO/2;  --SEGNALE A 0 PER MEZZO PERIODO
        CLOCK_50 <= '1';
        WAIT FOR PERIODO/2;  --SEGNALE A 1 PER MEZZO PERIODO
   END PROCESS;


   
   
END BEH;