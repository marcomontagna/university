
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_DLX_IR_SIZE32_PC_SIZE32 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_DLX_IR_SIZE32_PC_SIZE32;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_rbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_rbsh_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_rbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal MR_int_1_31_port, MR_int_1_30_port, MR_int_1_29_port, 
      MR_int_1_28_port, MR_int_1_27_port, MR_int_1_26_port, MR_int_1_25_port, 
      MR_int_1_24_port, MR_int_1_23_port, MR_int_1_22_port, MR_int_1_21_port, 
      MR_int_1_20_port, MR_int_1_19_port, MR_int_1_18_port, MR_int_1_17_port, 
      MR_int_1_16_port, MR_int_1_15_port, MR_int_1_14_port, MR_int_1_13_port, 
      MR_int_1_12_port, MR_int_1_11_port, MR_int_1_10_port, MR_int_1_9_port, 
      MR_int_1_8_port, MR_int_1_7_port, MR_int_1_6_port, MR_int_1_5_port, 
      MR_int_1_4_port, MR_int_1_3_port, MR_int_1_2_port, MR_int_1_1_port, 
      MR_int_1_0_port, MR_int_2_31_port, MR_int_2_30_port, MR_int_2_29_port, 
      MR_int_2_28_port, MR_int_2_27_port, MR_int_2_26_port, MR_int_2_25_port, 
      MR_int_2_24_port, MR_int_2_23_port, MR_int_2_22_port, MR_int_2_21_port, 
      MR_int_2_20_port, MR_int_2_19_port, MR_int_2_18_port, MR_int_2_17_port, 
      MR_int_2_16_port, MR_int_2_15_port, MR_int_2_14_port, MR_int_2_13_port, 
      MR_int_2_12_port, MR_int_2_11_port, MR_int_2_10_port, MR_int_2_9_port, 
      MR_int_2_8_port, MR_int_2_7_port, MR_int_2_6_port, MR_int_2_5_port, 
      MR_int_2_4_port, MR_int_2_3_port, MR_int_2_2_port, MR_int_2_1_port, 
      MR_int_2_0_port, MR_int_3_31_port, MR_int_3_30_port, MR_int_3_29_port, 
      MR_int_3_28_port, MR_int_3_27_port, MR_int_3_26_port, MR_int_3_25_port, 
      MR_int_3_24_port, MR_int_3_23_port, MR_int_3_22_port, MR_int_3_21_port, 
      MR_int_3_20_port, MR_int_3_19_port, MR_int_3_18_port, MR_int_3_17_port, 
      MR_int_3_16_port, MR_int_3_15_port, MR_int_3_14_port, MR_int_3_13_port, 
      MR_int_3_12_port, MR_int_3_11_port, MR_int_3_10_port, MR_int_3_9_port, 
      MR_int_3_8_port, MR_int_3_7_port, MR_int_3_6_port, MR_int_3_5_port, 
      MR_int_3_4_port, MR_int_3_3_port, MR_int_3_2_port, MR_int_3_1_port, 
      MR_int_3_0_port, MR_int_4_31_port, MR_int_4_30_port, MR_int_4_29_port, 
      MR_int_4_28_port, MR_int_4_27_port, MR_int_4_26_port, MR_int_4_25_port, 
      MR_int_4_24_port, MR_int_4_23_port, MR_int_4_22_port, MR_int_4_21_port, 
      MR_int_4_20_port, MR_int_4_19_port, MR_int_4_18_port, MR_int_4_17_port, 
      MR_int_4_16_port, MR_int_4_15_port, MR_int_4_14_port, MR_int_4_13_port, 
      MR_int_4_12_port, MR_int_4_11_port, MR_int_4_10_port, MR_int_4_9_port, 
      MR_int_4_8_port, MR_int_4_7_port, MR_int_4_6_port, MR_int_4_5_port, 
      MR_int_4_4_port, MR_int_4_3_port, MR_int_4_2_port, MR_int_4_1_port, 
      MR_int_4_0_port, n1, n2, n3 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => MR_int_4_31_port, B => MR_int_4_15_port, S 
                           => n3, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => MR_int_4_30_port, B => MR_int_4_14_port, S 
                           => n3, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => MR_int_4_29_port, B => MR_int_4_13_port, S 
                           => n3, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => MR_int_4_28_port, B => MR_int_4_12_port, S 
                           => n3, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => MR_int_4_27_port, B => MR_int_4_11_port, S 
                           => n3, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => MR_int_4_26_port, B => MR_int_4_10_port, S 
                           => n3, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => MR_int_4_25_port, B => MR_int_4_9_port, S 
                           => n3, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => MR_int_4_24_port, B => MR_int_4_8_port, S 
                           => n3, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => MR_int_4_23_port, B => MR_int_4_7_port, S 
                           => n2, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => MR_int_4_22_port, B => MR_int_4_6_port, S 
                           => n2, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => MR_int_4_21_port, B => MR_int_4_5_port, S 
                           => n2, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => MR_int_4_20_port, B => MR_int_4_4_port, S 
                           => n2, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => MR_int_4_19_port, B => MR_int_4_3_port, S 
                           => n2, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => MR_int_4_18_port, B => MR_int_4_2_port, S 
                           => n2, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => MR_int_4_17_port, B => MR_int_4_1_port, S 
                           => n2, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => MR_int_4_16_port, B => MR_int_4_0_port, S 
                           => n2, Z => B(16));
   M1_4_15 : MUX2_X1 port map( A => MR_int_4_15_port, B => MR_int_4_31_port, S 
                           => n2, Z => B(15));
   M1_4_14 : MUX2_X1 port map( A => MR_int_4_14_port, B => MR_int_4_30_port, S 
                           => n2, Z => B(14));
   M1_4_13 : MUX2_X1 port map( A => MR_int_4_13_port, B => MR_int_4_29_port, S 
                           => n2, Z => B(13));
   M1_4_12 : MUX2_X1 port map( A => MR_int_4_12_port, B => MR_int_4_28_port, S 
                           => n2, Z => B(12));
   M1_4_11 : MUX2_X1 port map( A => MR_int_4_11_port, B => MR_int_4_27_port, S 
                           => n1, Z => B(11));
   M1_4_10 : MUX2_X1 port map( A => MR_int_4_10_port, B => MR_int_4_26_port, S 
                           => n1, Z => B(10));
   M1_4_9 : MUX2_X1 port map( A => MR_int_4_9_port, B => MR_int_4_25_port, S =>
                           n1, Z => B(9));
   M1_4_8 : MUX2_X1 port map( A => MR_int_4_8_port, B => MR_int_4_24_port, S =>
                           n1, Z => B(8));
   M1_4_7 : MUX2_X1 port map( A => MR_int_4_7_port, B => MR_int_4_23_port, S =>
                           n1, Z => B(7));
   M1_4_6 : MUX2_X1 port map( A => MR_int_4_6_port, B => MR_int_4_22_port, S =>
                           n1, Z => B(6));
   M1_4_5 : MUX2_X1 port map( A => MR_int_4_5_port, B => MR_int_4_21_port, S =>
                           n1, Z => B(5));
   M1_4_4 : MUX2_X1 port map( A => MR_int_4_4_port, B => MR_int_4_20_port, S =>
                           n1, Z => B(4));
   M1_4_3 : MUX2_X1 port map( A => MR_int_4_3_port, B => MR_int_4_19_port, S =>
                           n1, Z => B(3));
   M1_4_2 : MUX2_X1 port map( A => MR_int_4_2_port, B => MR_int_4_18_port, S =>
                           n1, Z => B(2));
   M1_4_1 : MUX2_X1 port map( A => MR_int_4_1_port, B => MR_int_4_17_port, S =>
                           n1, Z => B(1));
   M1_4_0 : MUX2_X1 port map( A => MR_int_4_0_port, B => MR_int_4_16_port, S =>
                           n1, Z => B(0));
   M1_3_31_0 : MUX2_X1 port map( A => MR_int_3_31_port, B => MR_int_3_7_port, S
                           => SH(3), Z => MR_int_4_31_port);
   M1_3_30_0 : MUX2_X1 port map( A => MR_int_3_30_port, B => MR_int_3_6_port, S
                           => SH(3), Z => MR_int_4_30_port);
   M1_3_29_0 : MUX2_X1 port map( A => MR_int_3_29_port, B => MR_int_3_5_port, S
                           => SH(3), Z => MR_int_4_29_port);
   M1_3_28_0 : MUX2_X1 port map( A => MR_int_3_28_port, B => MR_int_3_4_port, S
                           => SH(3), Z => MR_int_4_28_port);
   M1_3_27_0 : MUX2_X1 port map( A => MR_int_3_27_port, B => MR_int_3_3_port, S
                           => SH(3), Z => MR_int_4_27_port);
   M1_3_26_0 : MUX2_X1 port map( A => MR_int_3_26_port, B => MR_int_3_2_port, S
                           => SH(3), Z => MR_int_4_26_port);
   M1_3_25_0 : MUX2_X1 port map( A => MR_int_3_25_port, B => MR_int_3_1_port, S
                           => SH(3), Z => MR_int_4_25_port);
   M1_3_24_0 : MUX2_X1 port map( A => MR_int_3_24_port, B => MR_int_3_0_port, S
                           => SH(3), Z => MR_int_4_24_port);
   M1_3_23_0 : MUX2_X1 port map( A => MR_int_3_23_port, B => MR_int_3_31_port, 
                           S => SH(3), Z => MR_int_4_23_port);
   M1_3_22_0 : MUX2_X1 port map( A => MR_int_3_22_port, B => MR_int_3_30_port, 
                           S => SH(3), Z => MR_int_4_22_port);
   M1_3_21_0 : MUX2_X1 port map( A => MR_int_3_21_port, B => MR_int_3_29_port, 
                           S => SH(3), Z => MR_int_4_21_port);
   M1_3_20_0 : MUX2_X1 port map( A => MR_int_3_20_port, B => MR_int_3_28_port, 
                           S => SH(3), Z => MR_int_4_20_port);
   M1_3_19_0 : MUX2_X1 port map( A => MR_int_3_19_port, B => MR_int_3_27_port, 
                           S => SH(3), Z => MR_int_4_19_port);
   M1_3_18_0 : MUX2_X1 port map( A => MR_int_3_18_port, B => MR_int_3_26_port, 
                           S => SH(3), Z => MR_int_4_18_port);
   M1_3_17_0 : MUX2_X1 port map( A => MR_int_3_17_port, B => MR_int_3_25_port, 
                           S => SH(3), Z => MR_int_4_17_port);
   M1_3_16_0 : MUX2_X1 port map( A => MR_int_3_16_port, B => MR_int_3_24_port, 
                           S => SH(3), Z => MR_int_4_16_port);
   M1_3_15_0 : MUX2_X1 port map( A => MR_int_3_15_port, B => MR_int_3_23_port, 
                           S => SH(3), Z => MR_int_4_15_port);
   M1_3_14_0 : MUX2_X1 port map( A => MR_int_3_14_port, B => MR_int_3_22_port, 
                           S => SH(3), Z => MR_int_4_14_port);
   M1_3_13_0 : MUX2_X1 port map( A => MR_int_3_13_port, B => MR_int_3_21_port, 
                           S => SH(3), Z => MR_int_4_13_port);
   M1_3_12_0 : MUX2_X1 port map( A => MR_int_3_12_port, B => MR_int_3_20_port, 
                           S => SH(3), Z => MR_int_4_12_port);
   M1_3_11_0 : MUX2_X1 port map( A => MR_int_3_11_port, B => MR_int_3_19_port, 
                           S => SH(3), Z => MR_int_4_11_port);
   M1_3_10_0 : MUX2_X1 port map( A => MR_int_3_10_port, B => MR_int_3_18_port, 
                           S => SH(3), Z => MR_int_4_10_port);
   M1_3_9_0 : MUX2_X1 port map( A => MR_int_3_9_port, B => MR_int_3_17_port, S 
                           => SH(3), Z => MR_int_4_9_port);
   M1_3_8_0 : MUX2_X1 port map( A => MR_int_3_8_port, B => MR_int_3_16_port, S 
                           => SH(3), Z => MR_int_4_8_port);
   M1_3_7 : MUX2_X1 port map( A => MR_int_3_7_port, B => MR_int_3_15_port, S =>
                           SH(3), Z => MR_int_4_7_port);
   M1_3_6 : MUX2_X1 port map( A => MR_int_3_6_port, B => MR_int_3_14_port, S =>
                           SH(3), Z => MR_int_4_6_port);
   M1_3_5 : MUX2_X1 port map( A => MR_int_3_5_port, B => MR_int_3_13_port, S =>
                           SH(3), Z => MR_int_4_5_port);
   M1_3_4 : MUX2_X1 port map( A => MR_int_3_4_port, B => MR_int_3_12_port, S =>
                           SH(3), Z => MR_int_4_4_port);
   M1_3_3 : MUX2_X1 port map( A => MR_int_3_3_port, B => MR_int_3_11_port, S =>
                           SH(3), Z => MR_int_4_3_port);
   M1_3_2 : MUX2_X1 port map( A => MR_int_3_2_port, B => MR_int_3_10_port, S =>
                           SH(3), Z => MR_int_4_2_port);
   M1_3_1 : MUX2_X1 port map( A => MR_int_3_1_port, B => MR_int_3_9_port, S => 
                           SH(3), Z => MR_int_4_1_port);
   M1_3_0 : MUX2_X1 port map( A => MR_int_3_0_port, B => MR_int_3_8_port, S => 
                           SH(3), Z => MR_int_4_0_port);
   M1_2_31_0 : MUX2_X1 port map( A => MR_int_2_31_port, B => MR_int_2_3_port, S
                           => SH(2), Z => MR_int_3_31_port);
   M1_2_30_0 : MUX2_X1 port map( A => MR_int_2_30_port, B => MR_int_2_2_port, S
                           => SH(2), Z => MR_int_3_30_port);
   M1_2_29_0 : MUX2_X1 port map( A => MR_int_2_29_port, B => MR_int_2_1_port, S
                           => SH(2), Z => MR_int_3_29_port);
   M1_2_28_0 : MUX2_X1 port map( A => MR_int_2_28_port, B => MR_int_2_0_port, S
                           => SH(2), Z => MR_int_3_28_port);
   M1_2_27_0 : MUX2_X1 port map( A => MR_int_2_27_port, B => MR_int_2_31_port, 
                           S => SH(2), Z => MR_int_3_27_port);
   M1_2_26_0 : MUX2_X1 port map( A => MR_int_2_26_port, B => MR_int_2_30_port, 
                           S => SH(2), Z => MR_int_3_26_port);
   M1_2_25_0 : MUX2_X1 port map( A => MR_int_2_25_port, B => MR_int_2_29_port, 
                           S => SH(2), Z => MR_int_3_25_port);
   M1_2_24_0 : MUX2_X1 port map( A => MR_int_2_24_port, B => MR_int_2_28_port, 
                           S => SH(2), Z => MR_int_3_24_port);
   M1_2_23_0 : MUX2_X1 port map( A => MR_int_2_23_port, B => MR_int_2_27_port, 
                           S => SH(2), Z => MR_int_3_23_port);
   M1_2_22_0 : MUX2_X1 port map( A => MR_int_2_22_port, B => MR_int_2_26_port, 
                           S => SH(2), Z => MR_int_3_22_port);
   M1_2_21_0 : MUX2_X1 port map( A => MR_int_2_21_port, B => MR_int_2_25_port, 
                           S => SH(2), Z => MR_int_3_21_port);
   M1_2_20_0 : MUX2_X1 port map( A => MR_int_2_20_port, B => MR_int_2_24_port, 
                           S => SH(2), Z => MR_int_3_20_port);
   M1_2_19_0 : MUX2_X1 port map( A => MR_int_2_19_port, B => MR_int_2_23_port, 
                           S => SH(2), Z => MR_int_3_19_port);
   M1_2_18_0 : MUX2_X1 port map( A => MR_int_2_18_port, B => MR_int_2_22_port, 
                           S => SH(2), Z => MR_int_3_18_port);
   M1_2_17_0 : MUX2_X1 port map( A => MR_int_2_17_port, B => MR_int_2_21_port, 
                           S => SH(2), Z => MR_int_3_17_port);
   M1_2_16_0 : MUX2_X1 port map( A => MR_int_2_16_port, B => MR_int_2_20_port, 
                           S => SH(2), Z => MR_int_3_16_port);
   M1_2_15_0 : MUX2_X1 port map( A => MR_int_2_15_port, B => MR_int_2_19_port, 
                           S => SH(2), Z => MR_int_3_15_port);
   M1_2_14_0 : MUX2_X1 port map( A => MR_int_2_14_port, B => MR_int_2_18_port, 
                           S => SH(2), Z => MR_int_3_14_port);
   M1_2_13_0 : MUX2_X1 port map( A => MR_int_2_13_port, B => MR_int_2_17_port, 
                           S => SH(2), Z => MR_int_3_13_port);
   M1_2_12_0 : MUX2_X1 port map( A => MR_int_2_12_port, B => MR_int_2_16_port, 
                           S => SH(2), Z => MR_int_3_12_port);
   M1_2_11_0 : MUX2_X1 port map( A => MR_int_2_11_port, B => MR_int_2_15_port, 
                           S => SH(2), Z => MR_int_3_11_port);
   M1_2_10_0 : MUX2_X1 port map( A => MR_int_2_10_port, B => MR_int_2_14_port, 
                           S => SH(2), Z => MR_int_3_10_port);
   M1_2_9_0 : MUX2_X1 port map( A => MR_int_2_9_port, B => MR_int_2_13_port, S 
                           => SH(2), Z => MR_int_3_9_port);
   M1_2_8_0 : MUX2_X1 port map( A => MR_int_2_8_port, B => MR_int_2_12_port, S 
                           => SH(2), Z => MR_int_3_8_port);
   M1_2_7_0 : MUX2_X1 port map( A => MR_int_2_7_port, B => MR_int_2_11_port, S 
                           => SH(2), Z => MR_int_3_7_port);
   M1_2_6_0 : MUX2_X1 port map( A => MR_int_2_6_port, B => MR_int_2_10_port, S 
                           => SH(2), Z => MR_int_3_6_port);
   M1_2_5_0 : MUX2_X1 port map( A => MR_int_2_5_port, B => MR_int_2_9_port, S 
                           => SH(2), Z => MR_int_3_5_port);
   M1_2_4_0 : MUX2_X1 port map( A => MR_int_2_4_port, B => MR_int_2_8_port, S 
                           => SH(2), Z => MR_int_3_4_port);
   M1_2_3 : MUX2_X1 port map( A => MR_int_2_3_port, B => MR_int_2_7_port, S => 
                           SH(2), Z => MR_int_3_3_port);
   M1_2_2 : MUX2_X1 port map( A => MR_int_2_2_port, B => MR_int_2_6_port, S => 
                           SH(2), Z => MR_int_3_2_port);
   M1_2_1 : MUX2_X1 port map( A => MR_int_2_1_port, B => MR_int_2_5_port, S => 
                           SH(2), Z => MR_int_3_1_port);
   M1_2_0 : MUX2_X1 port map( A => MR_int_2_0_port, B => MR_int_2_4_port, S => 
                           SH(2), Z => MR_int_3_0_port);
   M1_1_31_0 : MUX2_X1 port map( A => MR_int_1_31_port, B => MR_int_1_1_port, S
                           => SH(1), Z => MR_int_2_31_port);
   M1_1_30_0 : MUX2_X1 port map( A => MR_int_1_30_port, B => MR_int_1_0_port, S
                           => SH(1), Z => MR_int_2_30_port);
   M1_1_29_0 : MUX2_X1 port map( A => MR_int_1_29_port, B => MR_int_1_31_port, 
                           S => SH(1), Z => MR_int_2_29_port);
   M1_1_28_0 : MUX2_X1 port map( A => MR_int_1_28_port, B => MR_int_1_30_port, 
                           S => SH(1), Z => MR_int_2_28_port);
   M1_1_27_0 : MUX2_X1 port map( A => MR_int_1_27_port, B => MR_int_1_29_port, 
                           S => SH(1), Z => MR_int_2_27_port);
   M1_1_26_0 : MUX2_X1 port map( A => MR_int_1_26_port, B => MR_int_1_28_port, 
                           S => SH(1), Z => MR_int_2_26_port);
   M1_1_25_0 : MUX2_X1 port map( A => MR_int_1_25_port, B => MR_int_1_27_port, 
                           S => SH(1), Z => MR_int_2_25_port);
   M1_1_24_0 : MUX2_X1 port map( A => MR_int_1_24_port, B => MR_int_1_26_port, 
                           S => SH(1), Z => MR_int_2_24_port);
   M1_1_23_0 : MUX2_X1 port map( A => MR_int_1_23_port, B => MR_int_1_25_port, 
                           S => SH(1), Z => MR_int_2_23_port);
   M1_1_22_0 : MUX2_X1 port map( A => MR_int_1_22_port, B => MR_int_1_24_port, 
                           S => SH(1), Z => MR_int_2_22_port);
   M1_1_21_0 : MUX2_X1 port map( A => MR_int_1_21_port, B => MR_int_1_23_port, 
                           S => SH(1), Z => MR_int_2_21_port);
   M1_1_20_0 : MUX2_X1 port map( A => MR_int_1_20_port, B => MR_int_1_22_port, 
                           S => SH(1), Z => MR_int_2_20_port);
   M1_1_19_0 : MUX2_X1 port map( A => MR_int_1_19_port, B => MR_int_1_21_port, 
                           S => SH(1), Z => MR_int_2_19_port);
   M1_1_18_0 : MUX2_X1 port map( A => MR_int_1_18_port, B => MR_int_1_20_port, 
                           S => SH(1), Z => MR_int_2_18_port);
   M1_1_17_0 : MUX2_X1 port map( A => MR_int_1_17_port, B => MR_int_1_19_port, 
                           S => SH(1), Z => MR_int_2_17_port);
   M1_1_16_0 : MUX2_X1 port map( A => MR_int_1_16_port, B => MR_int_1_18_port, 
                           S => SH(1), Z => MR_int_2_16_port);
   M1_1_15_0 : MUX2_X1 port map( A => MR_int_1_15_port, B => MR_int_1_17_port, 
                           S => SH(1), Z => MR_int_2_15_port);
   M1_1_14_0 : MUX2_X1 port map( A => MR_int_1_14_port, B => MR_int_1_16_port, 
                           S => SH(1), Z => MR_int_2_14_port);
   M1_1_13_0 : MUX2_X1 port map( A => MR_int_1_13_port, B => MR_int_1_15_port, 
                           S => SH(1), Z => MR_int_2_13_port);
   M1_1_12_0 : MUX2_X1 port map( A => MR_int_1_12_port, B => MR_int_1_14_port, 
                           S => SH(1), Z => MR_int_2_12_port);
   M1_1_11_0 : MUX2_X1 port map( A => MR_int_1_11_port, B => MR_int_1_13_port, 
                           S => SH(1), Z => MR_int_2_11_port);
   M1_1_10_0 : MUX2_X1 port map( A => MR_int_1_10_port, B => MR_int_1_12_port, 
                           S => SH(1), Z => MR_int_2_10_port);
   M1_1_9_0 : MUX2_X1 port map( A => MR_int_1_9_port, B => MR_int_1_11_port, S 
                           => SH(1), Z => MR_int_2_9_port);
   M1_1_8_0 : MUX2_X1 port map( A => MR_int_1_8_port, B => MR_int_1_10_port, S 
                           => SH(1), Z => MR_int_2_8_port);
   M1_1_7_0 : MUX2_X1 port map( A => MR_int_1_7_port, B => MR_int_1_9_port, S 
                           => SH(1), Z => MR_int_2_7_port);
   M1_1_6_0 : MUX2_X1 port map( A => MR_int_1_6_port, B => MR_int_1_8_port, S 
                           => SH(1), Z => MR_int_2_6_port);
   M1_1_5_0 : MUX2_X1 port map( A => MR_int_1_5_port, B => MR_int_1_7_port, S 
                           => SH(1), Z => MR_int_2_5_port);
   M1_1_4_0 : MUX2_X1 port map( A => MR_int_1_4_port, B => MR_int_1_6_port, S 
                           => SH(1), Z => MR_int_2_4_port);
   M1_1_3_0 : MUX2_X1 port map( A => MR_int_1_3_port, B => MR_int_1_5_port, S 
                           => SH(1), Z => MR_int_2_3_port);
   M1_1_2_0 : MUX2_X1 port map( A => MR_int_1_2_port, B => MR_int_1_4_port, S 
                           => SH(1), Z => MR_int_2_2_port);
   M1_1_1 : MUX2_X1 port map( A => MR_int_1_1_port, B => MR_int_1_3_port, S => 
                           SH(1), Z => MR_int_2_1_port);
   M1_1_0 : MUX2_X1 port map( A => MR_int_1_0_port, B => MR_int_1_2_port, S => 
                           SH(1), Z => MR_int_2_0_port);
   M1_0_31_0 : MUX2_X1 port map( A => A(31), B => A(0), S => SH(0), Z => 
                           MR_int_1_31_port);
   M1_0_30_0 : MUX2_X1 port map( A => A(30), B => A(31), S => SH(0), Z => 
                           MR_int_1_30_port);
   M1_0_29_0 : MUX2_X1 port map( A => A(29), B => A(30), S => SH(0), Z => 
                           MR_int_1_29_port);
   M1_0_28_0 : MUX2_X1 port map( A => A(28), B => A(29), S => SH(0), Z => 
                           MR_int_1_28_port);
   M1_0_27_0 : MUX2_X1 port map( A => A(27), B => A(28), S => SH(0), Z => 
                           MR_int_1_27_port);
   M1_0_26_0 : MUX2_X1 port map( A => A(26), B => A(27), S => SH(0), Z => 
                           MR_int_1_26_port);
   M1_0_25_0 : MUX2_X1 port map( A => A(25), B => A(26), S => SH(0), Z => 
                           MR_int_1_25_port);
   M1_0_24_0 : MUX2_X1 port map( A => A(24), B => A(25), S => SH(0), Z => 
                           MR_int_1_24_port);
   M1_0_23_0 : MUX2_X1 port map( A => A(23), B => A(24), S => SH(0), Z => 
                           MR_int_1_23_port);
   M1_0_22_0 : MUX2_X1 port map( A => A(22), B => A(23), S => SH(0), Z => 
                           MR_int_1_22_port);
   M1_0_21_0 : MUX2_X1 port map( A => A(21), B => A(22), S => SH(0), Z => 
                           MR_int_1_21_port);
   M1_0_20_0 : MUX2_X1 port map( A => A(20), B => A(21), S => SH(0), Z => 
                           MR_int_1_20_port);
   M1_0_19_0 : MUX2_X1 port map( A => A(19), B => A(20), S => SH(0), Z => 
                           MR_int_1_19_port);
   M1_0_18_0 : MUX2_X1 port map( A => A(18), B => A(19), S => SH(0), Z => 
                           MR_int_1_18_port);
   M1_0_17_0 : MUX2_X1 port map( A => A(17), B => A(18), S => SH(0), Z => 
                           MR_int_1_17_port);
   M1_0_16_0 : MUX2_X1 port map( A => A(16), B => A(17), S => SH(0), Z => 
                           MR_int_1_16_port);
   M1_0_15_0 : MUX2_X1 port map( A => A(15), B => A(16), S => SH(0), Z => 
                           MR_int_1_15_port);
   M1_0_14_0 : MUX2_X1 port map( A => A(14), B => A(15), S => SH(0), Z => 
                           MR_int_1_14_port);
   M1_0_13_0 : MUX2_X1 port map( A => A(13), B => A(14), S => SH(0), Z => 
                           MR_int_1_13_port);
   M1_0_12_0 : MUX2_X1 port map( A => A(12), B => A(13), S => SH(0), Z => 
                           MR_int_1_12_port);
   M1_0_11_0 : MUX2_X1 port map( A => A(11), B => A(12), S => SH(0), Z => 
                           MR_int_1_11_port);
   M1_0_10_0 : MUX2_X1 port map( A => A(10), B => A(11), S => SH(0), Z => 
                           MR_int_1_10_port);
   M1_0_9_0 : MUX2_X1 port map( A => A(9), B => A(10), S => SH(0), Z => 
                           MR_int_1_9_port);
   M1_0_8_0 : MUX2_X1 port map( A => A(8), B => A(9), S => SH(0), Z => 
                           MR_int_1_8_port);
   M1_0_7_0 : MUX2_X1 port map( A => A(7), B => A(8), S => SH(0), Z => 
                           MR_int_1_7_port);
   M1_0_6_0 : MUX2_X1 port map( A => A(6), B => A(7), S => SH(0), Z => 
                           MR_int_1_6_port);
   M1_0_5_0 : MUX2_X1 port map( A => A(5), B => A(6), S => SH(0), Z => 
                           MR_int_1_5_port);
   M1_0_4_0 : MUX2_X1 port map( A => A(4), B => A(5), S => SH(0), Z => 
                           MR_int_1_4_port);
   M1_0_3_0 : MUX2_X1 port map( A => A(3), B => A(4), S => SH(0), Z => 
                           MR_int_1_3_port);
   M1_0_2_0 : MUX2_X1 port map( A => A(2), B => A(3), S => SH(0), Z => 
                           MR_int_1_2_port);
   M1_0_1_0 : MUX2_X1 port map( A => A(1), B => A(2), S => SH(0), Z => 
                           MR_int_1_1_port);
   M1_0_0 : MUX2_X1 port map( A => A(0), B => A(1), S => SH(0), Z => 
                           MR_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(4), Z => n1);
   U3 : BUF_X1 port map( A => SH(4), Z => n2);
   U4 : BUF_X1 port map( A => SH(4), Z => n3);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_lbsh_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_lbsh_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_lbsh_0 is

   component BUF_X1
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, 
      ML_int_1_28_port, ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, 
      ML_int_1_24_port, ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, 
      ML_int_1_20_port, ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, 
      ML_int_1_16_port, ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, 
      ML_int_1_12_port, ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, 
      ML_int_1_8_port, ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, 
      ML_int_1_4_port, ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, 
      ML_int_1_0_port, ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, 
      ML_int_2_28_port, ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, 
      ML_int_2_24_port, ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, 
      ML_int_2_20_port, ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, 
      ML_int_2_16_port, ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, 
      ML_int_2_12_port, ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, 
      ML_int_2_8_port, ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, 
      ML_int_2_4_port, ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, 
      ML_int_2_0_port, ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, 
      ML_int_3_28_port, ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, 
      ML_int_3_24_port, ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, 
      ML_int_3_20_port, ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, 
      ML_int_3_16_port, ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, 
      ML_int_3_12_port, ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, 
      ML_int_3_8_port, ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, 
      ML_int_3_4_port, ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, 
      ML_int_3_0_port, ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, 
      ML_int_4_28_port, ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, 
      ML_int_4_24_port, ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, 
      ML_int_4_20_port, ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, 
      ML_int_4_16_port, ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, 
      ML_int_4_12_port, ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, 
      ML_int_4_8_port, ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, 
      ML_int_4_4_port, ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, 
      ML_int_4_0_port, n1, n2, n3 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n3, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n3, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n3, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n3, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n3, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n3, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n3, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n3, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => n2, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => n2, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => n2, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => n2, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => n2, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => n2, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => n2, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => n2, Z => B(16));
   M0_4_15 : MUX2_X1 port map( A => ML_int_4_15_port, B => ML_int_4_31_port, S 
                           => n2, Z => B(15));
   M0_4_14 : MUX2_X1 port map( A => ML_int_4_14_port, B => ML_int_4_30_port, S 
                           => n2, Z => B(14));
   M0_4_13 : MUX2_X1 port map( A => ML_int_4_13_port, B => ML_int_4_29_port, S 
                           => n2, Z => B(13));
   M0_4_12 : MUX2_X1 port map( A => ML_int_4_12_port, B => ML_int_4_28_port, S 
                           => n2, Z => B(12));
   M0_4_11 : MUX2_X1 port map( A => ML_int_4_11_port, B => ML_int_4_27_port, S 
                           => n1, Z => B(11));
   M0_4_10 : MUX2_X1 port map( A => ML_int_4_10_port, B => ML_int_4_26_port, S 
                           => n1, Z => B(10));
   M0_4_9 : MUX2_X1 port map( A => ML_int_4_9_port, B => ML_int_4_25_port, S =>
                           n1, Z => B(9));
   M0_4_8 : MUX2_X1 port map( A => ML_int_4_8_port, B => ML_int_4_24_port, S =>
                           n1, Z => B(8));
   M0_4_7 : MUX2_X1 port map( A => ML_int_4_7_port, B => ML_int_4_23_port, S =>
                           n1, Z => B(7));
   M0_4_6 : MUX2_X1 port map( A => ML_int_4_6_port, B => ML_int_4_22_port, S =>
                           n1, Z => B(6));
   M0_4_5 : MUX2_X1 port map( A => ML_int_4_5_port, B => ML_int_4_21_port, S =>
                           n1, Z => B(5));
   M0_4_4 : MUX2_X1 port map( A => ML_int_4_4_port, B => ML_int_4_20_port, S =>
                           n1, Z => B(4));
   M0_4_3 : MUX2_X1 port map( A => ML_int_4_3_port, B => ML_int_4_19_port, S =>
                           n1, Z => B(3));
   M0_4_2 : MUX2_X1 port map( A => ML_int_4_2_port, B => ML_int_4_18_port, S =>
                           n1, Z => B(2));
   M0_4_1 : MUX2_X1 port map( A => ML_int_4_1_port, B => ML_int_4_17_port, S =>
                           n1, Z => B(1));
   M0_4_0 : MUX2_X1 port map( A => ML_int_4_0_port, B => ML_int_4_16_port, S =>
                           n1, Z => B(0));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => SH(3), Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => SH(3), Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => SH(3), Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => SH(3), Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => SH(3), Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => SH(3), Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => SH(3), Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => SH(3), Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => SH(3), Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => SH(3), Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => SH(3), Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => SH(3), Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => SH(3), Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => SH(3), Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => SH(3), Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => SH(3), Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => SH(3), Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => SH(3), Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => SH(3), Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => SH(3), Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => SH(3), Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => SH(3), Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           SH(3), Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           SH(3), Z => ML_int_4_8_port);
   M0_3_7 : MUX2_X1 port map( A => ML_int_3_7_port, B => ML_int_3_31_port, S =>
                           SH(3), Z => ML_int_4_7_port);
   M0_3_6 : MUX2_X1 port map( A => ML_int_3_6_port, B => ML_int_3_30_port, S =>
                           SH(3), Z => ML_int_4_6_port);
   M0_3_5 : MUX2_X1 port map( A => ML_int_3_5_port, B => ML_int_3_29_port, S =>
                           SH(3), Z => ML_int_4_5_port);
   M0_3_4 : MUX2_X1 port map( A => ML_int_3_4_port, B => ML_int_3_28_port, S =>
                           SH(3), Z => ML_int_4_4_port);
   M0_3_3 : MUX2_X1 port map( A => ML_int_3_3_port, B => ML_int_3_27_port, S =>
                           SH(3), Z => ML_int_4_3_port);
   M0_3_2 : MUX2_X1 port map( A => ML_int_3_2_port, B => ML_int_3_26_port, S =>
                           SH(3), Z => ML_int_4_2_port);
   M0_3_1 : MUX2_X1 port map( A => ML_int_3_1_port, B => ML_int_3_25_port, S =>
                           SH(3), Z => ML_int_4_1_port);
   M0_3_0 : MUX2_X1 port map( A => ML_int_3_0_port, B => ML_int_3_24_port, S =>
                           SH(3), Z => ML_int_4_0_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => SH(2), Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => SH(2), Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => SH(2), Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => SH(2), Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => SH(2), Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => SH(2), Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => SH(2), Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => SH(2), Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => SH(2), Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => SH(2), Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => SH(2), Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => SH(2), Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => SH(2), Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => SH(2), Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => SH(2), Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => SH(2), Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => SH(2), Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => SH(2), Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => SH(2), Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => SH(2), Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => SH(2), Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => SH(2), Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           SH(2), Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           SH(2), Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           SH(2), Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           SH(2), Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           SH(2), Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           SH(2), Z => ML_int_3_4_port);
   M0_2_3 : MUX2_X1 port map( A => ML_int_2_3_port, B => ML_int_2_31_port, S =>
                           SH(2), Z => ML_int_3_3_port);
   M0_2_2 : MUX2_X1 port map( A => ML_int_2_2_port, B => ML_int_2_30_port, S =>
                           SH(2), Z => ML_int_3_2_port);
   M0_2_1 : MUX2_X1 port map( A => ML_int_2_1_port, B => ML_int_2_29_port, S =>
                           SH(2), Z => ML_int_3_1_port);
   M0_2_0 : MUX2_X1 port map( A => ML_int_2_0_port, B => ML_int_2_28_port, S =>
                           SH(2), Z => ML_int_3_0_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => SH(1), Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => SH(1), Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => SH(1), Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => SH(1), Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => SH(1), Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => SH(1), Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => SH(1), Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => SH(1), Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => SH(1), Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => SH(1), Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => SH(1), Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => SH(1), Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => SH(1), Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => SH(1), Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => SH(1), Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => SH(1), Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => SH(1), Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => SH(1), Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => SH(1), Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => SH(1), Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => SH(1), Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => SH(1), Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           SH(1), Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           SH(1), Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           SH(1), Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           SH(1), Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           SH(1), Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           SH(1), Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           SH(1), Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           SH(1), Z => ML_int_2_2_port);
   M0_1_1 : MUX2_X1 port map( A => ML_int_1_1_port, B => ML_int_1_31_port, S =>
                           SH(1), Z => ML_int_2_1_port);
   M0_1_0 : MUX2_X1 port map( A => ML_int_1_0_port, B => ML_int_1_30_port, S =>
                           SH(1), Z => ML_int_2_0_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => SH(0), Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => SH(0), Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => SH(0), Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => SH(0), Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => SH(0), Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => SH(0), Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => SH(0), Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => SH(0), Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => SH(0), Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => SH(0), Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => SH(0), Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => SH(0), Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => SH(0), Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => SH(0), Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => SH(0), Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => SH(0), Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => SH(0), Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => SH(0), Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => SH(0), Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => SH(0), Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => SH(0), Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => SH(0), Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => SH(0), Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => SH(0), Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => SH(0), Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => SH(0), Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => SH(0), Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => SH(0), Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => SH(0), Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => SH(0), Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => SH(0), Z => 
                           ML_int_1_1_port);
   M0_0_0 : MUX2_X1 port map( A => A(0), B => A(31), S => SH(0), Z => 
                           ML_int_1_0_port);
   U2 : BUF_X1 port map( A => SH(4), Z => n1);
   U3 : BUF_X1 port map( A => SH(4), Z => n2);
   U4 : BUF_X1 port map( A => SH(4), Z => n3);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_sra_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_sra_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_sra_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, B_25_port, 
      B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, B_19_port, 
      B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, B_13_port, 
      B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port, B_6_port, 
      B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171 : std_logic;

begin
   B <= ( A(31), B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, B_0_port );
   
   U2 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n73);
   U3 : INV_X1 port map( A => SH(4), ZN => n1);
   U4 : OAI221_X1 port map( B1 => n2, B2 => n3, C1 => n4, C2 => n1, A => n5, ZN
                           => B_9_port);
   U5 : AOI222_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, C1 => n10, 
                           C2 => n11, ZN => n5);
   U6 : INV_X1 port map( A => n12, ZN => n2);
   U7 : OAI221_X1 port map( B1 => n13, B2 => n3, C1 => n14, C2 => n1, A => n15,
                           ZN => B_8_port);
   U8 : AOI222_X1 port map( A1 => n6, A2 => n16, B1 => n8, B2 => n17, C1 => n10
                           , C2 => n18, ZN => n15);
   U9 : INV_X1 port map( A => n19, ZN => n13);
   U10 : OAI221_X1 port map( B1 => n20, B2 => n3, C1 => n21, C2 => n1, A => n22
                           , ZN => B_7_port);
   U11 : AOI222_X1 port map( A1 => n6, A2 => n23, B1 => n8, B2 => n24, C1 => 
                           n10, C2 => n25, ZN => n22);
   U12 : OAI221_X1 port map( B1 => n26, B2 => n3, C1 => n27, C2 => n1, A => n28
                           , ZN => B_6_port);
   U13 : AOI222_X1 port map( A1 => n6, A2 => n29, B1 => n8, B2 => n30, C1 => 
                           n10, C2 => n31, ZN => n28);
   U14 : OAI221_X1 port map( B1 => n32, B2 => n3, C1 => n33, C2 => n1, A => n34
                           , ZN => B_5_port);
   U15 : AOI222_X1 port map( A1 => n6, A2 => n12, B1 => n8, B2 => n7, C1 => n10
                           , C2 => n9, ZN => n34);
   U16 : OAI221_X1 port map( B1 => n35, B2 => n3, C1 => n36, C2 => n1, A => n37
                           , ZN => B_4_port);
   U17 : AOI222_X1 port map( A1 => n6, A2 => n19, B1 => n8, B2 => n16, C1 => 
                           n10, C2 => n17, ZN => n37);
   U18 : OAI221_X1 port map( B1 => n20, B2 => n38, C1 => n39, C2 => n1, A => 
                           n40, ZN => B_3_port);
   U19 : AOI222_X1 port map( A1 => n10, A2 => n24, B1 => n41, B2 => n42, C1 => 
                           n8, C2 => n23, ZN => n40);
   U20 : OAI221_X1 port map( B1 => n43, B2 => n44, C1 => n45, C2 => n46, A => 
                           n47, ZN => n42);
   U21 : AOI22_X1 port map( A1 => A(5), A2 => n48, B1 => A(6), B2 => n49, ZN =>
                           n47);
   U22 : INV_X1 port map( A => A(4), ZN => n44);
   U23 : AOI221_X1 port map( B1 => n50, B2 => A(8), C1 => n51, C2 => A(7), A =>
                           n52, ZN => n20);
   U24 : OAI22_X1 port map( A1 => n53, A2 => n54, B1 => n55, B2 => n56, ZN => 
                           n52);
   U25 : OAI21_X1 port map( B1 => SH(4), B2 => n57, A => n58, ZN => B_30_port);
   U26 : OAI221_X1 port map( B1 => n26, B2 => n38, C1 => n59, C2 => n1, A => 
                           n60, ZN => B_2_port);
   U27 : AOI222_X1 port map( A1 => n10, A2 => n30, B1 => n41, B2 => n61, C1 => 
                           n8, C2 => n29, ZN => n60);
   U28 : OAI221_X1 port map( B1 => n43, B2 => n46, C1 => n45, C2 => n62, A => 
                           n63, ZN => n61);
   U29 : AOI22_X1 port map( A1 => A(4), A2 => n48, B1 => A(5), B2 => n49, ZN =>
                           n63);
   U30 : AOI221_X1 port map( B1 => n50, B2 => A(7), C1 => n51, C2 => A(6), A =>
                           n64, ZN => n26);
   U31 : OAI22_X1 port map( A1 => n65, A2 => n54, B1 => n53, B2 => n56, ZN => 
                           n64);
   U32 : OAI21_X1 port map( B1 => SH(4), B2 => n66, A => n58, ZN => B_29_port);
   U33 : OAI21_X1 port map( B1 => SH(4), B2 => n67, A => n58, ZN => B_28_port);
   U34 : OAI21_X1 port map( B1 => SH(4), B2 => n68, A => n58, ZN => B_27_port);
   U35 : OAI21_X1 port map( B1 => SH(4), B2 => n69, A => n58, ZN => B_26_port);
   U36 : OAI21_X1 port map( B1 => SH(4), B2 => n4, A => n58, ZN => B_25_port);
   U37 : AOI221_X1 port map( B1 => n70, B2 => n71, C1 => n72, C2 => n73, A => 
                           n74, ZN => n4);
   U38 : OAI21_X1 port map( B1 => SH(4), B2 => n14, A => n58, ZN => B_24_port);
   U39 : AOI221_X1 port map( B1 => n75, B2 => n71, C1 => n76, C2 => n73, A => 
                           n74, ZN => n14);
   U40 : OAI21_X1 port map( B1 => SH(4), B2 => n21, A => n58, ZN => B_23_port);
   U41 : AOI221_X1 port map( B1 => n77, B2 => n71, C1 => n78, C2 => n73, A => 
                           n74, ZN => n21);
   U42 : OAI21_X1 port map( B1 => SH(4), B2 => n27, A => n58, ZN => B_22_port);
   U43 : AOI221_X1 port map( B1 => n79, B2 => n71, C1 => n80, C2 => n73, A => 
                           n81, ZN => n27);
   U44 : INV_X1 port map( A => n82, ZN => n81);
   U45 : AOI21_X1 port map( B1 => n83, B2 => n84, A => n85, ZN => n82);
   U46 : OAI21_X1 port map( B1 => SH(4), B2 => n33, A => n58, ZN => B_21_port);
   U47 : AOI221_X1 port map( B1 => n72, B2 => n71, C1 => n11, C2 => n73, A => 
                           n86, ZN => n33);
   U48 : INV_X1 port map( A => n87, ZN => n86);
   U49 : AOI21_X1 port map( B1 => n83, B2 => n70, A => n85, ZN => n87);
   U50 : OAI21_X1 port map( B1 => SH(4), B2 => n36, A => n58, ZN => B_20_port);
   U51 : AOI221_X1 port map( B1 => n76, B2 => n71, C1 => n18, C2 => n73, A => 
                           n88, ZN => n36);
   U52 : INV_X1 port map( A => n89, ZN => n88);
   U53 : AOI21_X1 port map( B1 => n83, B2 => n75, A => n85, ZN => n89);
   U54 : OAI221_X1 port map( B1 => n32, B2 => n38, C1 => n90, C2 => n1, A => 
                           n91, ZN => B_1_port);
   U55 : AOI222_X1 port map( A1 => n10, A2 => n7, B1 => n41, B2 => n92, C1 => 
                           n8, C2 => n12, ZN => n91);
   U56 : OAI221_X1 port map( B1 => n43, B2 => n55, C1 => n45, C2 => n53, A => 
                           n93, ZN => n12);
   U57 : AOI22_X1 port map( A1 => A(11), A2 => n48, B1 => A(12), B2 => n49, ZN 
                           => n93);
   U58 : OAI221_X1 port map( B1 => n43, B2 => n62, C1 => n45, C2 => n94, A => 
                           n95, ZN => n92);
   U59 : AOI22_X1 port map( A1 => A(3), A2 => n48, B1 => A(4), B2 => n49, ZN =>
                           n95);
   U60 : INV_X1 port map( A => A(1), ZN => n94);
   U61 : AOI221_X1 port map( B1 => n50, B2 => A(6), C1 => n51, C2 => A(5), A =>
                           n96, ZN => n32);
   U62 : OAI22_X1 port map( A1 => n97, A2 => n54, B1 => n65, B2 => n56, ZN => 
                           n96);
   U63 : OAI21_X1 port map( B1 => SH(4), B2 => n39, A => n58, ZN => B_19_port);
   U64 : AOI221_X1 port map( B1 => n78, B2 => n71, C1 => n25, C2 => n73, A => 
                           n98, ZN => n39);
   U65 : INV_X1 port map( A => n99, ZN => n98);
   U66 : AOI21_X1 port map( B1 => n83, B2 => n77, A => n85, ZN => n99);
   U67 : NOR2_X1 port map( A1 => n100, A2 => n101, ZN => n85);
   U68 : OAI21_X1 port map( B1 => SH(4), B2 => n59, A => n58, ZN => B_18_port);
   U69 : AOI221_X1 port map( B1 => n80, B2 => n71, C1 => n31, C2 => n73, A => 
                           n102, ZN => n59);
   U70 : INV_X1 port map( A => n103, ZN => n102);
   U71 : AOI22_X1 port map( A1 => n104, A2 => n84, B1 => n83, B2 => n79, ZN => 
                           n103);
   U72 : OAI21_X1 port map( B1 => SH(4), B2 => n90, A => n58, ZN => B_17_port);
   U73 : AOI221_X1 port map( B1 => n11, B2 => n71, C1 => n9, C2 => n73, A => 
                           n105, ZN => n90);
   U74 : INV_X1 port map( A => n106, ZN => n105);
   U75 : AOI22_X1 port map( A1 => n104, A2 => n70, B1 => n83, B2 => n72, ZN => 
                           n106);
   U76 : OAI21_X1 port map( B1 => SH(4), B2 => n107, A => n58, ZN => B_16_port)
                           ;
   U77 : OAI221_X1 port map( B1 => n108, B2 => n38, C1 => n109, C2 => n3, A => 
                           n110, ZN => B_15_port);
   U78 : AOI221_X1 port map( B1 => n10, B2 => n77, C1 => n8, C2 => n78, A => 
                           n111, ZN => n110);
   U79 : INV_X1 port map( A => n58, ZN => n111);
   U80 : NAND2_X1 port map( A1 => SH(4), A2 => A(31), ZN => n58);
   U81 : INV_X1 port map( A => n25, ZN => n108);
   U82 : OAI221_X1 port map( B1 => n112, B2 => n3, C1 => n57, C2 => n1, A => 
                           n113, ZN => B_14_port);
   U83 : AOI222_X1 port map( A1 => n6, A2 => n31, B1 => n8, B2 => n80, C1 => 
                           n10, C2 => n79, ZN => n113);
   U84 : AOI21_X1 port map( B1 => n84, B2 => n73, A => n114, ZN => n57);
   U85 : OAI221_X1 port map( B1 => n115, B2 => n3, C1 => n66, C2 => n1, A => 
                           n116, ZN => B_13_port);
   U86 : AOI222_X1 port map( A1 => n6, A2 => n9, B1 => n8, B2 => n11, C1 => n10
                           , C2 => n72, ZN => n116);
   U87 : OAI221_X1 port map( B1 => n43, B2 => n117, C1 => n45, C2 => n118, A =>
                           n119, ZN => n72);
   U88 : AOI22_X1 port map( A1 => A(27), A2 => n48, B1 => A(28), B2 => n49, ZN 
                           => n119);
   U89 : OAI221_X1 port map( B1 => n43, B2 => n120, C1 => n45, C2 => n121, A =>
                           n122, ZN => n11);
   U90 : AOI22_X1 port map( A1 => A(23), A2 => n48, B1 => A(24), B2 => n49, ZN 
                           => n122);
   U91 : OAI221_X1 port map( B1 => n43, B2 => n123, C1 => n45, C2 => n124, A =>
                           n125, ZN => n9);
   U92 : AOI22_X1 port map( A1 => A(19), A2 => n48, B1 => A(20), B2 => n49, ZN 
                           => n125);
   U93 : AOI21_X1 port map( B1 => n70, B2 => n73, A => n114, ZN => n66);
   U94 : INV_X1 port map( A => n126, ZN => n70);
   U95 : AOI222_X1 port map( A1 => n51, A2 => A(29), B1 => n50, B2 => A(30), C1
                           => SH(1), C2 => A(31), ZN => n126);
   U96 : INV_X1 port map( A => n7, ZN => n115);
   U97 : OAI221_X1 port map( B1 => n43, B2 => n127, C1 => n45, C2 => n128, A =>
                           n129, ZN => n7);
   U98 : AOI22_X1 port map( A1 => A(15), A2 => n48, B1 => A(16), B2 => n49, ZN 
                           => n129);
   U99 : INV_X1 port map( A => A(14), ZN => n127);
   U100 : OAI221_X1 port map( B1 => n130, B2 => n3, C1 => n67, C2 => n1, A => 
                           n131, ZN => B_12_port);
   U101 : AOI222_X1 port map( A1 => n6, A2 => n17, B1 => n8, B2 => n18, C1 => 
                           n10, C2 => n76, ZN => n131);
   U102 : AOI21_X1 port map( B1 => n75, B2 => n73, A => n114, ZN => n67);
   U103 : INV_X1 port map( A => n16, ZN => n130);
   U104 : OAI221_X1 port map( B1 => n132, B2 => n3, C1 => n68, C2 => n1, A => 
                           n133, ZN => B_11_port);
   U105 : AOI222_X1 port map( A1 => n6, A2 => n24, B1 => n8, B2 => n25, C1 => 
                           n10, C2 => n78, ZN => n133);
   U106 : OAI221_X1 port map( B1 => n43, B2 => n134, C1 => n45, C2 => n135, A 
                           => n136, ZN => n78);
   U107 : AOI22_X1 port map( A1 => A(25), A2 => n48, B1 => A(26), B2 => n49, ZN
                           => n136);
   U108 : OAI221_X1 port map( B1 => n137, B2 => n43, C1 => n138, C2 => n45, A 
                           => n139, ZN => n25);
   U109 : AOI22_X1 port map( A1 => A(21), A2 => n48, B1 => A(22), B2 => n49, ZN
                           => n139);
   U110 : INV_X1 port map( A => n109, ZN => n24);
   U111 : AOI221_X1 port map( B1 => n50, B2 => A(16), C1 => n51, C2 => A(15), A
                           => n140, ZN => n109);
   U112 : OAI22_X1 port map( A1 => n124, A2 => n54, B1 => n123, B2 => n56, ZN 
                           => n140);
   U113 : INV_X1 port map( A => A(17), ZN => n124);
   U114 : AOI21_X1 port map( B1 => n77, B2 => n73, A => n114, ZN => n68);
   U115 : OAI21_X1 port map( B1 => n101, B2 => n141, A => n100, ZN => n114);
   U116 : INV_X1 port map( A => A(31), ZN => n141);
   U117 : OAI221_X1 port map( B1 => n43, B2 => n142, C1 => n45, C2 => n143, A 
                           => n144, ZN => n77);
   U118 : AOI22_X1 port map( A1 => A(29), A2 => n48, B1 => A(30), B2 => n49, ZN
                           => n144);
   U119 : INV_X1 port map( A => n23, ZN => n132);
   U120 : OAI221_X1 port map( B1 => n43, B2 => n145, C1 => n45, C2 => n146, A 
                           => n147, ZN => n23);
   U121 : AOI22_X1 port map( A1 => A(13), A2 => n48, B1 => A(14), B2 => n49, ZN
                           => n147);
   U122 : OAI221_X1 port map( B1 => n148, B2 => n3, C1 => n69, C2 => n1, A => 
                           n149, ZN => B_10_port);
   U123 : AOI222_X1 port map( A1 => n6, A2 => n30, B1 => n8, B2 => n31, C1 => 
                           n10, C2 => n80, ZN => n149);
   U124 : OAI221_X1 port map( B1 => n43, B2 => n135, C1 => n45, C2 => n120, A 
                           => n150, ZN => n80);
   U125 : AOI22_X1 port map( A1 => A(24), A2 => n48, B1 => A(25), B2 => n49, ZN
                           => n150);
   U126 : INV_X1 port map( A => A(22), ZN => n120);
   U127 : INV_X1 port map( A => A(23), ZN => n135);
   U128 : OAI221_X1 port map( B1 => n138, B2 => n43, C1 => n123, C2 => n45, A 
                           => n151, ZN => n31);
   U129 : AOI22_X1 port map( A1 => A(20), A2 => n48, B1 => A(21), B2 => n49, ZN
                           => n151);
   U130 : INV_X1 port map( A => n112, ZN => n30);
   U131 : AOI221_X1 port map( B1 => n50, B2 => A(15), C1 => n51, C2 => A(14), A
                           => n152, ZN => n112);
   U132 : INV_X1 port map( A => n153, ZN => n152);
   U133 : AOI22_X1 port map( A1 => A(16), A2 => n48, B1 => A(17), B2 => n49, ZN
                           => n153);
   U134 : INV_X1 port map( A => n38, ZN => n6);
   U135 : AOI221_X1 port map( B1 => n84, B2 => n71, C1 => n79, C2 => n73, A => 
                           n74, ZN => n69);
   U136 : INV_X1 port map( A => n100, ZN => n74);
   U137 : NAND2_X1 port map( A1 => A(31), A2 => SH(3), ZN => n100);
   U138 : OAI221_X1 port map( B1 => n43, B2 => n143, C1 => n45, C2 => n117, A 
                           => n154, ZN => n79);
   U139 : AOI22_X1 port map( A1 => A(28), A2 => n48, B1 => A(29), B2 => n49, ZN
                           => n154);
   U140 : INV_X1 port map( A => A(26), ZN => n117);
   U141 : INV_X1 port map( A => A(27), ZN => n143);
   U142 : MUX2_X1 port map( A => A(31), B => A(30), S => n51, Z => n84);
   U143 : INV_X1 port map( A => n29, ZN => n148);
   U144 : OAI221_X1 port map( B1 => n43, B2 => n146, C1 => n45, C2 => n55, A =>
                           n155, ZN => n29);
   U145 : AOI22_X1 port map( A1 => A(12), A2 => n48, B1 => A(13), B2 => n49, ZN
                           => n155);
   U146 : INV_X1 port map( A => A(10), ZN => n55);
   U147 : INV_X1 port map( A => A(11), ZN => n146);
   U148 : OAI221_X1 port map( B1 => n35, B2 => n38, C1 => n107, C2 => n1, A => 
                           n156, ZN => B_0_port);
   U149 : AOI222_X1 port map( A1 => n10, A2 => n16, B1 => n41, B2 => n157, C1 
                           => n8, C2 => n19, ZN => n156);
   U150 : OAI221_X1 port map( B1 => n43, B2 => n53, C1 => n45, C2 => n65, A => 
                           n158, ZN => n19);
   U151 : AOI22_X1 port map( A1 => A(10), A2 => n48, B1 => A(11), B2 => n49, ZN
                           => n158);
   U152 : INV_X1 port map( A => A(8), ZN => n65);
   U153 : INV_X1 port map( A => A(9), ZN => n53);
   U154 : AND2_X1 port map( A1 => n159, A2 => n101, ZN => n8);
   U155 : OAI221_X1 port map( B1 => n54, B2 => n62, C1 => n56, C2 => n46, A => 
                           n160, ZN => n157);
   U156 : AOI22_X1 port map( A1 => A(1), A2 => n50, B1 => A(0), B2 => n51, ZN 
                           => n160);
   U157 : INV_X1 port map( A => A(3), ZN => n46);
   U158 : INV_X1 port map( A => A(2), ZN => n62);
   U159 : INV_X1 port map( A => n3, ZN => n41);
   U160 : NAND2_X1 port map( A1 => n73, A2 => n1, ZN => n3);
   U161 : OAI221_X1 port map( B1 => n43, B2 => n128, C1 => n45, C2 => n145, A 
                           => n161, ZN => n16);
   U162 : AOI22_X1 port map( A1 => A(14), A2 => n48, B1 => A(15), B2 => n49, ZN
                           => n161);
   U163 : INV_X1 port map( A => A(12), ZN => n145);
   U164 : INV_X1 port map( A => A(13), ZN => n128);
   U165 : AND2_X1 port map( A1 => SH(2), A2 => n159, ZN => n10);
   U166 : AND2_X1 port map( A1 => SH(3), A2 => n1, ZN => n159);
   U167 : AOI221_X1 port map( B1 => n18, B2 => n71, C1 => n17, C2 => n73, A => 
                           n162, ZN => n107);
   U168 : INV_X1 port map( A => n163, ZN => n162);
   U169 : AOI22_X1 port map( A1 => n104, A2 => n75, B1 => n83, B2 => n76, ZN =>
                           n163);
   U170 : OAI221_X1 port map( B1 => n43, B2 => n118, C1 => n45, C2 => n134, A 
                           => n164, ZN => n76);
   U171 : AOI22_X1 port map( A1 => A(26), A2 => n48, B1 => A(27), B2 => n49, ZN
                           => n164);
   U172 : INV_X1 port map( A => A(24), ZN => n134);
   U173 : INV_X1 port map( A => A(25), ZN => n118);
   U174 : AND2_X1 port map( A1 => SH(3), A2 => n101, ZN => n83);
   U175 : OAI221_X1 port map( B1 => n43, B2 => n165, C1 => n45, C2 => n142, A 
                           => n166, ZN => n75);
   U176 : AOI22_X1 port map( A1 => A(30), A2 => n48, B1 => A(31), B2 => n49, ZN
                           => n166);
   U177 : INV_X1 port map( A => A(28), ZN => n142);
   U178 : INV_X1 port map( A => A(29), ZN => n165);
   U179 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n104);
   U180 : OAI221_X1 port map( B1 => n54, B2 => n123, C1 => n138, C2 => n56, A 
                           => n167, ZN => n17);
   U181 : AOI22_X1 port map( A1 => A(17), A2 => n50, B1 => A(16), B2 => n51, ZN
                           => n167);
   U182 : INV_X1 port map( A => A(19), ZN => n138);
   U183 : INV_X1 port map( A => A(18), ZN => n123);
   U184 : OAI221_X1 port map( B1 => n43, B2 => n121, C1 => n137, C2 => n45, A 
                           => n168, ZN => n18);
   U185 : AOI22_X1 port map( A1 => A(22), A2 => n48, B1 => A(23), B2 => n49, ZN
                           => n168);
   U186 : INV_X1 port map( A => n56, ZN => n49);
   U187 : INV_X1 port map( A => n54, ZN => n48);
   U188 : INV_X1 port map( A => n51, ZN => n45);
   U189 : INV_X1 port map( A => A(20), ZN => n137);
   U190 : INV_X1 port map( A => A(21), ZN => n121);
   U191 : INV_X1 port map( A => n50, ZN => n43);
   U192 : NAND2_X1 port map( A1 => n71, A2 => n1, ZN => n38);
   U193 : NOR2_X1 port map( A1 => n101, A2 => SH(3), ZN => n71);
   U194 : INV_X1 port map( A => SH(2), ZN => n101);
   U195 : AOI221_X1 port map( B1 => n50, B2 => A(5), C1 => n51, C2 => A(4), A 
                           => n169, ZN => n35);
   U196 : OAI22_X1 port map( A1 => n170, A2 => n54, B1 => n97, B2 => n56, ZN =>
                           n169);
   U197 : NAND2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n56);
   U198 : INV_X1 port map( A => A(7), ZN => n97);
   U199 : NAND2_X1 port map( A1 => SH(1), A2 => n171, ZN => n54);
   U200 : INV_X1 port map( A => A(6), ZN => n170);
   U201 : NOR2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n51);
   U202 : NOR2_X1 port map( A1 => n171, A2 => SH(1), ZN => n50);
   U203 : INV_X1 port map( A => SH(0), ZN => n171);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_rash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32_DW_rash_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_rash_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, 
      n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, 
      n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, 
      n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, 
      n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, 
      n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, 
      n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162 : 
      std_logic;

begin
   
   U3 : NOR2_X2 port map( A1 => SH(0), A2 => SH(1), ZN => n50);
   U4 : NOR2_X2 port map( A1 => n162, A2 => SH(1), ZN => n49);
   U5 : INV_X1 port map( A => SH(4), ZN => n1);
   U6 : OAI221_X1 port map( B1 => n2, B2 => n3, C1 => n4, C2 => n1, A => n5, ZN
                           => B(9));
   U7 : AOI222_X1 port map( A1 => n6, A2 => n7, B1 => n8, B2 => n9, C1 => n10, 
                           C2 => n11, ZN => n5);
   U8 : OAI221_X1 port map( B1 => n12, B2 => n3, C1 => n13, C2 => n1, A => n14,
                           ZN => B(8));
   U9 : AOI222_X1 port map( A1 => n6, A2 => n15, B1 => n8, B2 => n16, C1 => n10
                           , C2 => n17, ZN => n14);
   U10 : OAI221_X1 port map( B1 => n18, B2 => n3, C1 => n19, C2 => n1, A => n20
                           , ZN => B(7));
   U11 : AOI222_X1 port map( A1 => n6, A2 => n21, B1 => n8, B2 => n22, C1 => 
                           n10, C2 => n23, ZN => n20);
   U12 : OAI221_X1 port map( B1 => n24, B2 => n3, C1 => n25, C2 => n1, A => n26
                           , ZN => B(6));
   U13 : AOI222_X1 port map( A1 => n6, A2 => n27, B1 => n8, B2 => n28, C1 => 
                           n10, C2 => n29, ZN => n26);
   U14 : OAI221_X1 port map( B1 => n30, B2 => n3, C1 => n31, C2 => n1, A => n32
                           , ZN => B(5));
   U15 : AOI222_X1 port map( A1 => n6, A2 => n33, B1 => n8, B2 => n7, C1 => n10
                           , C2 => n9, ZN => n32);
   U16 : OAI221_X1 port map( B1 => n34, B2 => n3, C1 => n35, C2 => n1, A => n36
                           , ZN => B(4));
   U17 : AOI222_X1 port map( A1 => n6, A2 => n37, B1 => n8, B2 => n15, C1 => 
                           n10, C2 => n16, ZN => n36);
   U18 : OAI221_X1 port map( B1 => n18, B2 => n38, C1 => n39, C2 => n1, A => 
                           n40, ZN => B(3));
   U19 : AOI222_X1 port map( A1 => n10, A2 => n22, B1 => n41, B2 => n42, C1 => 
                           n8, C2 => n21, ZN => n40);
   U20 : INV_X1 port map( A => n43, ZN => n21);
   U21 : OAI221_X1 port map( B1 => n44, B2 => n45, C1 => n46, C2 => n47, A => 
                           n48, ZN => n42);
   U22 : AOI22_X1 port map( A1 => A(4), A2 => n49, B1 => A(3), B2 => n50, ZN =>
                           n48);
   U23 : AOI221_X1 port map( B1 => n51, B2 => A(10), C1 => n52, C2 => A(9), A 
                           => n53, ZN => n18);
   U24 : OAI22_X1 port map( A1 => n54, A2 => n55, B1 => n56, B2 => n57, ZN => 
                           n53);
   U25 : AND2_X1 port map( A1 => n41, A2 => n58, ZN => B(31));
   U26 : AND2_X1 port map( A1 => n59, A2 => n41, ZN => B(30));
   U27 : OAI221_X1 port map( B1 => n24, B2 => n38, C1 => n60, C2 => n1, A => 
                           n61, ZN => B(2));
   U28 : AOI222_X1 port map( A1 => n10, A2 => n28, B1 => n41, B2 => n62, C1 => 
                           n8, C2 => n27, ZN => n61);
   U29 : INV_X1 port map( A => n63, ZN => n27);
   U30 : OAI221_X1 port map( B1 => n44, B2 => n47, C1 => n46, C2 => n64, A => 
                           n65, ZN => n62);
   U31 : AOI22_X1 port map( A1 => A(3), A2 => n49, B1 => A(2), B2 => n50, ZN =>
                           n65);
   U32 : AOI221_X1 port map( B1 => n51, B2 => A(9), C1 => n52, C2 => A(8), A =>
                           n66, ZN => n24);
   U33 : OAI22_X1 port map( A1 => n56, A2 => n55, B1 => n45, B2 => n57, ZN => 
                           n66);
   U34 : INV_X1 port map( A => A(7), ZN => n56);
   U35 : AND2_X1 port map( A1 => n67, A2 => n41, ZN => B(29));
   U36 : AND2_X1 port map( A1 => n68, A2 => n41, ZN => B(28));
   U37 : NOR3_X1 port map( A1 => n69, A2 => SH(4), A3 => SH(3), ZN => B(27));
   U38 : NOR2_X1 port map( A1 => SH(4), A2 => n70, ZN => B(26));
   U39 : NOR2_X1 port map( A1 => SH(4), A2 => n4, ZN => B(25));
   U40 : AOI22_X1 port map( A1 => n71, A2 => n72, B1 => n67, B2 => n73, ZN => 
                           n4);
   U41 : NOR2_X1 port map( A1 => SH(4), A2 => n13, ZN => B(24));
   U42 : AOI22_X1 port map( A1 => n74, A2 => n72, B1 => n68, B2 => n73, ZN => 
                           n13);
   U43 : NOR2_X1 port map( A1 => SH(4), A2 => n19, ZN => B(23));
   U44 : AOI222_X1 port map( A1 => n75, A2 => n73, B1 => n58, B2 => n76, C1 => 
                           n77, C2 => n72, ZN => n19);
   U45 : NOR2_X1 port map( A1 => SH(4), A2 => n25, ZN => B(22));
   U46 : AOI222_X1 port map( A1 => n78, A2 => n73, B1 => n59, B2 => n76, C1 => 
                           n79, C2 => n72, ZN => n25);
   U47 : NOR2_X1 port map( A1 => SH(4), A2 => n31, ZN => B(21));
   U48 : AOI222_X1 port map( A1 => n71, A2 => n73, B1 => n67, B2 => n76, C1 => 
                           n11, C2 => n72, ZN => n31);
   U49 : NOR2_X1 port map( A1 => SH(4), A2 => n35, ZN => B(20));
   U50 : AOI222_X1 port map( A1 => n74, A2 => n73, B1 => n68, B2 => n76, C1 => 
                           n17, C2 => n72, ZN => n35);
   U51 : OAI221_X1 port map( B1 => n30, B2 => n38, C1 => n80, C2 => n1, A => 
                           n81, ZN => B(1));
   U52 : AOI222_X1 port map( A1 => n10, A2 => n7, B1 => n41, B2 => n82, C1 => 
                           n8, C2 => n33, ZN => n81);
   U53 : INV_X1 port map( A => n2, ZN => n33);
   U54 : AOI221_X1 port map( B1 => n51, B2 => A(12), C1 => n52, C2 => A(11), A 
                           => n83, ZN => n2);
   U55 : OAI22_X1 port map( A1 => n84, A2 => n55, B1 => n85, B2 => n57, ZN => 
                           n83);
   U56 : OAI221_X1 port map( B1 => n44, B2 => n64, C1 => n46, C2 => n86, A => 
                           n87, ZN => n82);
   U57 : AOI22_X1 port map( A1 => A(2), A2 => n49, B1 => A(1), B2 => n50, ZN =>
                           n87);
   U58 : AOI221_X1 port map( B1 => n51, B2 => A(8), C1 => n52, C2 => A(7), A =>
                           n88, ZN => n30);
   U59 : OAI22_X1 port map( A1 => n45, A2 => n55, B1 => n47, B2 => n57, ZN => 
                           n88);
   U60 : INV_X1 port map( A => A(6), ZN => n45);
   U61 : NOR2_X1 port map( A1 => SH(4), A2 => n39, ZN => B(19));
   U62 : AOI222_X1 port map( A1 => n23, A2 => n72, B1 => n77, B2 => n73, C1 => 
                           n89, C2 => SH(3), ZN => n39);
   U63 : NOR2_X1 port map( A1 => SH(4), A2 => n60, ZN => B(18));
   U64 : AOI221_X1 port map( B1 => n79, B2 => n73, C1 => n29, C2 => n72, A => 
                           n90, ZN => n60);
   U65 : INV_X1 port map( A => n91, ZN => n90);
   U66 : AOI22_X1 port map( A1 => n92, A2 => n59, B1 => n76, B2 => n78, ZN => 
                           n91);
   U67 : NOR2_X1 port map( A1 => SH(4), A2 => n80, ZN => B(17));
   U68 : AOI221_X1 port map( B1 => n11, B2 => n73, C1 => n9, C2 => n72, A => 
                           n93, ZN => n80);
   U69 : INV_X1 port map( A => n94, ZN => n93);
   U70 : AOI22_X1 port map( A1 => n92, A2 => n67, B1 => n76, B2 => n71, ZN => 
                           n94);
   U71 : NOR2_X1 port map( A1 => SH(4), A2 => n95, ZN => B(16));
   U72 : OAI221_X1 port map( B1 => n96, B2 => n38, C1 => n97, C2 => n3, A => 
                           n98, ZN => B(15));
   U73 : AOI222_X1 port map( A1 => n10, A2 => n75, B1 => n99, B2 => n58, C1 => 
                           n8, C2 => n77, ZN => n98);
   U74 : INV_X1 port map( A => n23, ZN => n96);
   U75 : OAI221_X1 port map( B1 => n100, B2 => n38, C1 => n101, C2 => n3, A => 
                           n102, ZN => B(14));
   U76 : AOI222_X1 port map( A1 => n10, A2 => n78, B1 => n99, B2 => n59, C1 => 
                           n8, C2 => n79, ZN => n102);
   U77 : INV_X1 port map( A => n28, ZN => n101);
   U78 : INV_X1 port map( A => n29, ZN => n100);
   U79 : OAI221_X1 port map( B1 => n103, B2 => n38, C1 => n104, C2 => n3, A => 
                           n105, ZN => B(13));
   U80 : AOI222_X1 port map( A1 => n10, A2 => n71, B1 => n99, B2 => n67, C1 => 
                           n8, C2 => n11, ZN => n105);
   U81 : OAI221_X1 port map( B1 => n44, B2 => n106, C1 => n46, C2 => n107, A =>
                           n108, ZN => n11);
   U82 : AOI22_X1 port map( A1 => A(22), A2 => n49, B1 => A(21), B2 => n50, ZN 
                           => n108);
   U83 : INV_X1 port map( A => A(23), ZN => n107);
   U84 : OAI222_X1 port map( A1 => n55, A2 => n109, B1 => n46, B2 => n110, C1 
                           => n57, C2 => n111, ZN => n67);
   U85 : OAI221_X1 port map( B1 => n44, B2 => n112, C1 => n46, C2 => n113, A =>
                           n114, ZN => n71);
   U86 : AOI22_X1 port map( A1 => A(26), A2 => n49, B1 => A(25), B2 => n50, ZN 
                           => n114);
   U87 : INV_X1 port map( A => n7, ZN => n104);
   U88 : OAI221_X1 port map( B1 => n44, B2 => n115, C1 => n46, C2 => n116, A =>
                           n117, ZN => n7);
   U89 : AOI22_X1 port map( A1 => A(14), A2 => n49, B1 => A(13), B2 => n50, ZN 
                           => n117);
   U90 : INV_X1 port map( A => n9, ZN => n103);
   U91 : OAI221_X1 port map( B1 => n44, B2 => n118, C1 => n46, C2 => n119, A =>
                           n120, ZN => n9);
   U92 : AOI22_X1 port map( A1 => A(18), A2 => n49, B1 => A(17), B2 => n50, ZN 
                           => n120);
   U93 : INV_X1 port map( A => n121, ZN => B(12));
   U94 : AOI221_X1 port map( B1 => n16, B2 => n6, C1 => n15, C2 => n41, A => 
                           n122, ZN => n121);
   U95 : INV_X1 port map( A => n123, ZN => n122);
   U96 : AOI222_X1 port map( A1 => n10, A2 => n74, B1 => n99, B2 => n68, C1 => 
                           n8, C2 => n17, ZN => n123);
   U97 : NOR2_X1 port map( A1 => n1, A2 => n124, ZN => n99);
   U98 : OAI221_X1 port map( B1 => n97, B2 => n38, C1 => n43, C2 => n3, A => 
                           n125, ZN => B(11));
   U99 : AOI221_X1 port map( B1 => n10, B2 => n77, C1 => n8, C2 => n23, A => 
                           n126, ZN => n125);
   U100 : NOR3_X1 port map( A1 => n1, A2 => SH(3), A3 => n69, ZN => n126);
   U101 : INV_X1 port map( A => n89, ZN => n69);
   U102 : MUX2_X1 port map( A => n75, B => n58, S => SH(2), Z => n89);
   U103 : NOR2_X1 port map( A1 => n110, A2 => n57, ZN => n58);
   U104 : OAI221_X1 port map( B1 => n44, B2 => n109, C1 => n46, C2 => n111, A 
                           => n127, ZN => n75);
   U105 : AOI22_X1 port map( A1 => A(28), A2 => n49, B1 => A(27), B2 => n50, ZN
                           => n127);
   U106 : OAI221_X1 port map( B1 => n118, B2 => n55, C1 => n119, C2 => n57, A 
                           => n128, ZN => n23);
   U107 : AOI22_X1 port map( A1 => A(22), A2 => n51, B1 => A(21), B2 => n52, ZN
                           => n128);
   U108 : OAI221_X1 port map( B1 => n44, B2 => n129, C1 => n46, C2 => n130, A 
                           => n131, ZN => n77);
   U109 : AOI22_X1 port map( A1 => A(24), A2 => n49, B1 => A(23), B2 => n50, ZN
                           => n131);
   U110 : AOI221_X1 port map( B1 => n51, B2 => A(14), C1 => n52, C2 => A(13), A
                           => n132, ZN => n43);
   U111 : OAI22_X1 port map( A1 => n133, A2 => n55, B1 => n134, B2 => n57, ZN 
                           => n132);
   U112 : INV_X1 port map( A => A(12), ZN => n133);
   U113 : INV_X1 port map( A => n22, ZN => n97);
   U114 : OAI221_X1 port map( B1 => n44, B2 => n135, C1 => n46, C2 => n136, A 
                           => n137, ZN => n22);
   U115 : AOI22_X1 port map( A1 => A(16), A2 => n49, B1 => A(15), B2 => n50, ZN
                           => n137);
   U116 : OAI221_X1 port map( B1 => n63, B2 => n3, C1 => n70, C2 => n1, A => 
                           n138, ZN => B(10));
   U117 : AOI222_X1 port map( A1 => n6, A2 => n28, B1 => n8, B2 => n29, C1 => 
                           n10, C2 => n79, ZN => n138);
   U118 : OAI221_X1 port map( B1 => n44, B2 => n130, C1 => n46, C2 => n106, A 
                           => n139, ZN => n79);
   U119 : AOI22_X1 port map( A1 => A(23), A2 => n49, B1 => A(22), B2 => n50, ZN
                           => n139);
   U120 : INV_X1 port map( A => A(24), ZN => n106);
   U121 : INV_X1 port map( A => A(25), ZN => n130);
   U122 : OAI221_X1 port map( B1 => n119, B2 => n55, C1 => n135, C2 => n57, A 
                           => n140, ZN => n29);
   U123 : AOI22_X1 port map( A1 => A(21), A2 => n51, B1 => n52, B2 => A(20), ZN
                           => n140);
   U124 : OAI221_X1 port map( B1 => n44, B2 => n136, C1 => n46, C2 => n115, A 
                           => n141, ZN => n28);
   U125 : AOI22_X1 port map( A1 => A(15), A2 => n49, B1 => A(14), B2 => n50, ZN
                           => n141);
   U126 : INV_X1 port map( A => A(16), ZN => n115);
   U127 : INV_X1 port map( A => A(17), ZN => n136);
   U128 : INV_X1 port map( A => n38, ZN => n6);
   U129 : AOI22_X1 port map( A1 => n78, A2 => n72, B1 => n59, B2 => n73, ZN => 
                           n70);
   U130 : OAI22_X1 port map( A1 => n57, A2 => n109, B1 => n55, B2 => n110, ZN 
                           => n59);
   U131 : OAI221_X1 port map( B1 => n44, B2 => n111, C1 => n46, C2 => n112, A 
                           => n142, ZN => n78);
   U132 : AOI22_X1 port map( A1 => A(27), A2 => n49, B1 => A(26), B2 => n50, ZN
                           => n142);
   U133 : INV_X1 port map( A => A(28), ZN => n112);
   U134 : INV_X1 port map( A => A(29), ZN => n111);
   U135 : AOI221_X1 port map( B1 => n51, B2 => A(13), C1 => n52, C2 => A(12), A
                           => n143, ZN => n63);
   U136 : OAI22_X1 port map( A1 => n134, A2 => n55, B1 => n84, B2 => n57, ZN =>
                           n143);
   U137 : INV_X1 port map( A => A(10), ZN => n84);
   U138 : INV_X1 port map( A => A(11), ZN => n134);
   U139 : OAI221_X1 port map( B1 => n34, B2 => n38, C1 => n95, C2 => n1, A => 
                           n144, ZN => B(0));
   U140 : AOI222_X1 port map( A1 => n10, A2 => n15, B1 => n41, B2 => n145, C1 
                           => n8, C2 => n37, ZN => n144);
   U141 : INV_X1 port map( A => n12, ZN => n37);
   U142 : AOI221_X1 port map( B1 => n51, B2 => A(11), C1 => n52, C2 => A(10), A
                           => n146, ZN => n12);
   U143 : OAI22_X1 port map( A1 => n85, A2 => n55, B1 => n54, B2 => n57, ZN => 
                           n146);
   U144 : INV_X1 port map( A => A(8), ZN => n54);
   U145 : INV_X1 port map( A => A(9), ZN => n85);
   U146 : AND2_X1 port map( A1 => n147, A2 => n148, ZN => n8);
   U147 : OAI221_X1 port map( B1 => n44, B2 => n86, C1 => n46, C2 => n149, A =>
                           n150, ZN => n145);
   U148 : AOI22_X1 port map( A1 => A(1), A2 => n49, B1 => A(0), B2 => n50, ZN 
                           => n150);
   U149 : INV_X1 port map( A => A(2), ZN => n149);
   U150 : INV_X1 port map( A => A(3), ZN => n86);
   U151 : INV_X1 port map( A => n3, ZN => n41);
   U152 : NAND2_X1 port map( A1 => n72, A2 => n1, ZN => n3);
   U153 : OAI221_X1 port map( B1 => n44, B2 => n116, C1 => n46, C2 => n151, A 
                           => n152, ZN => n15);
   U154 : AOI22_X1 port map( A1 => A(13), A2 => n49, B1 => A(12), B2 => n50, ZN
                           => n152);
   U155 : INV_X1 port map( A => A(14), ZN => n151);
   U156 : INV_X1 port map( A => A(15), ZN => n116);
   U157 : AND2_X1 port map( A1 => SH(2), A2 => n147, ZN => n10);
   U158 : NOR2_X1 port map( A1 => n153, A2 => SH(4), ZN => n147);
   U159 : AOI221_X1 port map( B1 => n17, B2 => n73, C1 => n16, C2 => n72, A => 
                           n154, ZN => n95);
   U160 : INV_X1 port map( A => n155, ZN => n154);
   U161 : AOI22_X1 port map( A1 => n92, A2 => n68, B1 => n76, B2 => n74, ZN => 
                           n155);
   U162 : OAI221_X1 port map( B1 => n44, B2 => n113, C1 => n46, C2 => n129, A 
                           => n156, ZN => n74);
   U163 : AOI22_X1 port map( A1 => A(25), A2 => n49, B1 => A(24), B2 => n50, ZN
                           => n156);
   U164 : INV_X1 port map( A => A(26), ZN => n129);
   U165 : INV_X1 port map( A => A(27), ZN => n113);
   U166 : NOR2_X1 port map( A1 => n153, A2 => SH(2), ZN => n76);
   U167 : OAI221_X1 port map( B1 => n44, B2 => n110, C1 => n46, C2 => n109, A 
                           => n157, ZN => n68);
   U168 : AOI22_X1 port map( A1 => A(29), A2 => n49, B1 => A(28), B2 => n50, ZN
                           => n157);
   U169 : INV_X1 port map( A => A(30), ZN => n109);
   U170 : INV_X1 port map( A => A(31), ZN => n110);
   U171 : NOR2_X1 port map( A1 => n148, A2 => n153, ZN => n92);
   U172 : INV_X1 port map( A => n124, ZN => n72);
   U173 : NAND2_X1 port map( A1 => n148, A2 => n153, ZN => n124);
   U174 : INV_X1 port map( A => SH(3), ZN => n153);
   U175 : OAI221_X1 port map( B1 => n44, B2 => n119, C1 => n46, C2 => n135, A 
                           => n158, ZN => n16);
   U176 : AOI22_X1 port map( A1 => A(17), A2 => n49, B1 => A(16), B2 => n50, ZN
                           => n158);
   U177 : INV_X1 port map( A => A(18), ZN => n135);
   U178 : INV_X1 port map( A => A(19), ZN => n119);
   U179 : OAI221_X1 port map( B1 => n55, B2 => n159, C1 => n118, C2 => n57, A 
                           => n160, ZN => n17);
   U180 : AOI22_X1 port map( A1 => A(23), A2 => n51, B1 => A(22), B2 => n52, ZN
                           => n160);
   U181 : INV_X1 port map( A => A(20), ZN => n118);
   U182 : INV_X1 port map( A => A(21), ZN => n159);
   U183 : NAND2_X1 port map( A1 => n73, A2 => n1, ZN => n38);
   U184 : NOR2_X1 port map( A1 => n148, A2 => SH(3), ZN => n73);
   U185 : INV_X1 port map( A => SH(2), ZN => n148);
   U186 : AOI221_X1 port map( B1 => n51, B2 => A(7), C1 => n52, C2 => A(6), A 
                           => n161, ZN => n34);
   U187 : OAI22_X1 port map( A1 => n47, A2 => n55, B1 => n64, B2 => n57, ZN => 
                           n161);
   U188 : INV_X1 port map( A => n50, ZN => n57);
   U189 : INV_X1 port map( A => A(4), ZN => n64);
   U190 : INV_X1 port map( A => n49, ZN => n55);
   U191 : INV_X1 port map( A => A(5), ZN => n47);
   U192 : INV_X1 port map( A => n46, ZN => n52);
   U193 : NAND2_X1 port map( A1 => SH(1), A2 => n162, ZN => n46);
   U194 : INV_X1 port map( A => SH(0), ZN => n162);
   U195 : INV_X1 port map( A => n44, ZN => n51);
   U196 : NAND2_X1 port map( A1 => SH(1), A2 => SH(0), ZN => n44);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW_sla_0 is

   port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4 
         downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 downto
         0));

end SHIFTER_GENERIC_N32_DW_sla_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW_sla_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, n1, n2, n3, 
      n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
      n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34
      , n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, 
      n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63
      , n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, 
      n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92
      , n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, 
      n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, 
      n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, 
      n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, 
      n142, n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, 
      n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, 
      n166, n167, n168, n169, n170, n171, n172, n173 : std_logic;

begin
   B <= ( B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, B_26_port, 
      B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, B_20_port, 
      B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, B_14_port, 
      B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port, B_7_port,
      B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, A(0) );
   
   U2 : NOR2_X2 port map( A1 => SH(2), A2 => SH(3), ZN => n75);
   U3 : INV_X1 port map( A => SH(4), ZN => n1);
   U4 : OAI21_X1 port map( B1 => SH(4), B2 => n2, A => n3, ZN => B_9_port);
   U5 : OAI21_X1 port map( B1 => SH(4), B2 => n4, A => n3, ZN => B_8_port);
   U6 : OAI21_X1 port map( B1 => SH(4), B2 => n5, A => n3, ZN => B_7_port);
   U7 : OAI21_X1 port map( B1 => SH(4), B2 => n6, A => n3, ZN => B_6_port);
   U8 : OAI21_X1 port map( B1 => SH(4), B2 => n7, A => n3, ZN => B_5_port);
   U9 : OAI21_X1 port map( B1 => SH(4), B2 => n8, A => n3, ZN => B_4_port);
   U10 : OAI21_X1 port map( B1 => SH(4), B2 => n9, A => n3, ZN => B_3_port);
   U11 : OAI221_X1 port map( B1 => n10, B2 => n11, C1 => n12, C2 => n1, A => 
                           n13, ZN => B_31_port);
   U12 : AOI222_X1 port map( A1 => n14, A2 => n15, B1 => n16, B2 => n17, C1 => 
                           n18, C2 => n19, ZN => n13);
   U13 : OAI221_X1 port map( B1 => n20, B2 => n21, C1 => n22, C2 => n23, A => 
                           n24, ZN => n17);
   U14 : AOI22_X1 port map( A1 => A(30), A2 => n25, B1 => A(31), B2 => n26, ZN 
                           => n24);
   U15 : OAI221_X1 port map( B1 => n27, B2 => n11, C1 => n28, C2 => n1, A => 
                           n29, ZN => B_30_port);
   U16 : AOI222_X1 port map( A1 => n14, A2 => n30, B1 => n16, B2 => n31, C1 => 
                           n18, C2 => n32, ZN => n29);
   U17 : OAI221_X1 port map( B1 => n33, B2 => n21, C1 => n34, C2 => n35, A => 
                           n36, ZN => n31);
   U18 : AOI22_X1 port map( A1 => A(28), A2 => n37, B1 => A(27), B2 => n38, ZN 
                           => n36);
   U19 : INV_X1 port map( A => A(30), ZN => n35);
   U20 : OAI21_X1 port map( B1 => SH(4), B2 => n39, A => n3, ZN => B_2_port);
   U21 : OAI221_X1 port map( B1 => n40, B2 => n11, C1 => n41, C2 => n1, A => 
                           n42, ZN => B_29_port);
   U22 : AOI222_X1 port map( A1 => n14, A2 => n43, B1 => n16, B2 => n44, C1 => 
                           n18, C2 => n45, ZN => n42);
   U23 : OAI221_X1 port map( B1 => n33, B2 => n23, C1 => n34, C2 => n21, A => 
                           n46, ZN => n44);
   U24 : AOI22_X1 port map( A1 => A(27), A2 => n37, B1 => A(26), B2 => n38, ZN 
                           => n46);
   U25 : INV_X1 port map( A => A(29), ZN => n21);
   U26 : OAI221_X1 port map( B1 => n47, B2 => n11, C1 => n48, C2 => n1, A => 
                           n49, ZN => B_28_port);
   U27 : AOI222_X1 port map( A1 => n14, A2 => n50, B1 => n16, B2 => n51, C1 => 
                           n18, C2 => n52, ZN => n49);
   U28 : OAI221_X1 port map( B1 => n33, B2 => n53, C1 => n34, C2 => n23, A => 
                           n54, ZN => n51);
   U29 : AOI22_X1 port map( A1 => A(26), A2 => n37, B1 => A(25), B2 => n38, ZN 
                           => n54);
   U30 : INV_X1 port map( A => A(28), ZN => n23);
   U31 : INV_X1 port map( A => A(27), ZN => n53);
   U32 : INV_X1 port map( A => n55, ZN => n16);
   U33 : OAI221_X1 port map( B1 => n10, B2 => n55, C1 => n56, C2 => n1, A => 
                           n57, ZN => B_27_port);
   U34 : AOI222_X1 port map( A1 => n58, A2 => n19, B1 => n18, B2 => n15, C1 => 
                           n14, C2 => n59, ZN => n57);
   U35 : INV_X1 port map( A => n60, ZN => n19);
   U36 : AOI221_X1 port map( B1 => n25, B2 => A(26), C1 => n26, C2 => A(27), A 
                           => n61, ZN => n10);
   U37 : INV_X1 port map( A => n62, ZN => n61);
   U38 : AOI22_X1 port map( A1 => A(25), A2 => n37, B1 => A(24), B2 => n38, ZN 
                           => n62);
   U39 : OAI221_X1 port map( B1 => n27, B2 => n55, C1 => n63, C2 => n1, A => 
                           n64, ZN => B_26_port);
   U40 : AOI222_X1 port map( A1 => n58, A2 => n32, B1 => n18, B2 => n30, C1 => 
                           n14, C2 => n65, ZN => n64);
   U41 : INV_X1 port map( A => n66, ZN => n32);
   U42 : AOI221_X1 port map( B1 => n25, B2 => A(25), C1 => n26, C2 => A(26), A 
                           => n67, ZN => n27);
   U43 : INV_X1 port map( A => n68, ZN => n67);
   U44 : AOI22_X1 port map( A1 => A(24), A2 => n37, B1 => A(23), B2 => n38, ZN 
                           => n68);
   U45 : OAI221_X1 port map( B1 => n40, B2 => n55, C1 => n2, C2 => n1, A => n69
                           , ZN => B_25_port);
   U46 : AOI222_X1 port map( A1 => n58, A2 => n45, B1 => n18, B2 => n43, C1 => 
                           n14, C2 => n70, ZN => n69);
   U47 : INV_X1 port map( A => n71, ZN => n45);
   U48 : AOI221_X1 port map( B1 => n72, B2 => n73, C1 => n74, C2 => n75, A => 
                           n76, ZN => n2);
   U49 : INV_X1 port map( A => n77, ZN => n76);
   U50 : AOI21_X1 port map( B1 => n78, B2 => n79, A => n80, ZN => n77);
   U51 : AOI221_X1 port map( B1 => n25, B2 => A(24), C1 => n26, C2 => A(25), A 
                           => n81, ZN => n40);
   U52 : INV_X1 port map( A => n82, ZN => n81);
   U53 : AOI22_X1 port map( A1 => A(23), A2 => n37, B1 => A(22), B2 => n38, ZN 
                           => n82);
   U54 : OAI221_X1 port map( B1 => n47, B2 => n55, C1 => n4, C2 => n1, A => n83
                           , ZN => B_24_port);
   U55 : AOI222_X1 port map( A1 => n58, A2 => n52, B1 => n18, B2 => n50, C1 => 
                           n14, C2 => n84, ZN => n83);
   U56 : INV_X1 port map( A => n85, ZN => n52);
   U57 : AOI221_X1 port map( B1 => n86, B2 => n73, C1 => n87, C2 => n75, A => 
                           n88, ZN => n4);
   U58 : AOI221_X1 port map( B1 => n25, B2 => A(23), C1 => n26, C2 => A(24), A 
                           => n89, ZN => n47);
   U59 : INV_X1 port map( A => n90, ZN => n89);
   U60 : AOI22_X1 port map( A1 => A(22), A2 => n37, B1 => A(21), B2 => n38, ZN 
                           => n90);
   U61 : OAI221_X1 port map( B1 => n60, B2 => n55, C1 => n5, C2 => n1, A => n91
                           , ZN => B_23_port);
   U62 : AOI222_X1 port map( A1 => n58, A2 => n15, B1 => n18, B2 => n59, C1 => 
                           n14, C2 => n92, ZN => n91);
   U63 : INV_X1 port map( A => n93, ZN => n15);
   U64 : AOI221_X1 port map( B1 => n94, B2 => n73, C1 => n95, C2 => n75, A => 
                           n88, ZN => n5);
   U65 : AOI221_X1 port map( B1 => n25, B2 => A(22), C1 => n26, C2 => A(23), A 
                           => n96, ZN => n60);
   U66 : INV_X1 port map( A => n97, ZN => n96);
   U67 : AOI22_X1 port map( A1 => A(21), A2 => n37, B1 => A(20), B2 => n38, ZN 
                           => n97);
   U68 : OAI221_X1 port map( B1 => n66, B2 => n55, C1 => n6, C2 => n1, A => n98
                           , ZN => B_22_port);
   U69 : AOI222_X1 port map( A1 => n58, A2 => n30, B1 => n18, B2 => n65, C1 => 
                           n14, C2 => n99, ZN => n98);
   U70 : INV_X1 port map( A => n100, ZN => n30);
   U71 : AOI221_X1 port map( B1 => n101, B2 => n73, C1 => n102, C2 => n75, A =>
                           n88, ZN => n6);
   U72 : AOI221_X1 port map( B1 => n25, B2 => A(21), C1 => n26, C2 => A(22), A 
                           => n103, ZN => n66);
   U73 : INV_X1 port map( A => n104, ZN => n103);
   U74 : AOI22_X1 port map( A1 => A(20), A2 => n37, B1 => A(19), B2 => n38, ZN 
                           => n104);
   U75 : OAI221_X1 port map( B1 => n71, B2 => n55, C1 => n7, C2 => n1, A => 
                           n105, ZN => B_21_port);
   U76 : AOI222_X1 port map( A1 => n58, A2 => n43, B1 => n18, B2 => n70, C1 => 
                           n14, C2 => n74, ZN => n105);
   U77 : INV_X1 port map( A => n106, ZN => n43);
   U78 : AOI221_X1 port map( B1 => n79, B2 => n73, C1 => n72, C2 => n75, A => 
                           n88, ZN => n7);
   U79 : INV_X1 port map( A => n107, ZN => n88);
   U80 : AOI221_X1 port map( B1 => n25, B2 => A(20), C1 => n26, C2 => A(21), A 
                           => n108, ZN => n71);
   U81 : OAI22_X1 port map( A1 => n109, A2 => n20, B1 => n110, B2 => n22, ZN =>
                           n108);
   U82 : INV_X1 port map( A => A(19), ZN => n109);
   U83 : OAI221_X1 port map( B1 => n85, B2 => n55, C1 => n8, C2 => n1, A => 
                           n111, ZN => B_20_port);
   U84 : AOI222_X1 port map( A1 => n58, A2 => n50, B1 => n18, B2 => n84, C1 => 
                           n14, C2 => n87, ZN => n111);
   U85 : INV_X1 port map( A => n112, ZN => n50);
   U86 : AOI21_X1 port map( B1 => n86, B2 => n75, A => n113, ZN => n8);
   U87 : AOI221_X1 port map( B1 => n25, B2 => A(19), C1 => n26, C2 => A(20), A 
                           => n114, ZN => n85);
   U88 : OAI22_X1 port map( A1 => n110, A2 => n20, B1 => n115, B2 => n22, ZN =>
                           n114);
   U89 : INV_X1 port map( A => A(18), ZN => n110);
   U90 : OAI21_X1 port map( B1 => SH(4), B2 => n116, A => n3, ZN => B_1_port);
   U91 : OAI221_X1 port map( B1 => n93, B2 => n55, C1 => n9, C2 => n1, A => 
                           n117, ZN => B_19_port);
   U92 : AOI222_X1 port map( A1 => n58, A2 => n59, B1 => n18, B2 => n92, C1 => 
                           n14, C2 => n95, ZN => n117);
   U93 : AOI21_X1 port map( B1 => n94, B2 => n75, A => n113, ZN => n9);
   U94 : AOI221_X1 port map( B1 => n25, B2 => A(18), C1 => n26, C2 => A(19), A 
                           => n118, ZN => n93);
   U95 : OAI22_X1 port map( A1 => n115, A2 => n20, B1 => n119, B2 => n22, ZN =>
                           n118);
   U96 : INV_X1 port map( A => A(17), ZN => n115);
   U97 : OAI221_X1 port map( B1 => n100, B2 => n55, C1 => n39, C2 => n1, A => 
                           n120, ZN => B_18_port);
   U98 : AOI222_X1 port map( A1 => n58, A2 => n65, B1 => n18, B2 => n99, C1 => 
                           n14, C2 => n102, ZN => n120);
   U99 : AOI21_X1 port map( B1 => n101, B2 => n75, A => n113, ZN => n39);
   U100 : AOI221_X1 port map( B1 => n25, B2 => A(17), C1 => n26, C2 => A(18), A
                           => n121, ZN => n100);
   U101 : OAI22_X1 port map( A1 => n119, A2 => n20, B1 => n122, B2 => n22, ZN 
                           => n121);
   U102 : INV_X1 port map( A => A(16), ZN => n119);
   U103 : OAI221_X1 port map( B1 => n106, B2 => n55, C1 => n116, C2 => n1, A =>
                           n123, ZN => B_17_port);
   U104 : AOI222_X1 port map( A1 => n58, A2 => n70, B1 => n18, B2 => n74, C1 =>
                           n14, C2 => n72, ZN => n123);
   U105 : INV_X1 port map( A => n11, ZN => n58);
   U106 : AOI21_X1 port map( B1 => n79, B2 => n75, A => n113, ZN => n116);
   U107 : OAI21_X1 port map( B1 => n124, B2 => n125, A => n107, ZN => n113);
   U108 : AOI221_X1 port map( B1 => n25, B2 => A(16), C1 => n26, C2 => A(17), A
                           => n126, ZN => n106);
   U109 : OAI22_X1 port map( A1 => n122, A2 => n20, B1 => n127, B2 => n22, ZN 
                           => n126);
   U110 : OAI221_X1 port map( B1 => n128, B2 => n11, C1 => n112, C2 => n55, A 
                           => n129, ZN => B_16_port);
   U111 : AOI221_X1 port map( B1 => n14, B2 => n86, C1 => n18, C2 => n87, A => 
                           n130, ZN => n129);
   U112 : INV_X1 port map( A => n3, ZN => n130);
   U113 : AND2_X1 port map( A1 => n131, A2 => n125, ZN => n18);
   U114 : AND2_X1 port map( A1 => n131, A2 => SH(2), ZN => n14);
   U115 : AND2_X1 port map( A1 => SH(3), A2 => n1, ZN => n131);
   U116 : NAND2_X1 port map( A1 => n75, A2 => n1, ZN => n55);
   U117 : AOI221_X1 port map( B1 => n25, B2 => A(15), C1 => n26, C2 => A(16), A
                           => n132, ZN => n112);
   U118 : OAI22_X1 port map( A1 => n127, A2 => n20, B1 => n133, B2 => n22, ZN 
                           => n132);
   U119 : NAND2_X1 port map( A1 => n73, A2 => n1, ZN => n11);
   U120 : INV_X1 port map( A => n84, ZN => n128);
   U121 : OAI21_X1 port map( B1 => SH(4), B2 => n12, A => n3, ZN => B_15_port);
   U122 : AOI221_X1 port map( B1 => n92, B2 => n73, C1 => n59, C2 => n75, A => 
                           n134, ZN => n12);
   U123 : INV_X1 port map( A => n135, ZN => n134);
   U124 : AOI22_X1 port map( A1 => n136, A2 => n94, B1 => n78, B2 => n95, ZN =>
                           n135);
   U125 : OAI221_X1 port map( B1 => n33, B2 => n127, C1 => n34, C2 => n122, A 
                           => n137, ZN => n59);
   U126 : AOI22_X1 port map( A1 => A(13), A2 => n37, B1 => A(12), B2 => n38, ZN
                           => n137);
   U127 : INV_X1 port map( A => A(15), ZN => n122);
   U128 : OAI21_X1 port map( B1 => SH(4), B2 => n28, A => n3, ZN => B_14_port);
   U129 : AOI221_X1 port map( B1 => n99, B2 => n73, C1 => n65, C2 => n75, A => 
                           n138, ZN => n28);
   U130 : INV_X1 port map( A => n139, ZN => n138);
   U131 : AOI22_X1 port map( A1 => n136, A2 => n101, B1 => n78, B2 => n102, ZN 
                           => n139);
   U132 : OAI221_X1 port map( B1 => n33, B2 => n133, C1 => n34, C2 => n127, A 
                           => n140, ZN => n65);
   U133 : AOI22_X1 port map( A1 => A(12), A2 => n37, B1 => A(11), B2 => n38, ZN
                           => n140);
   U134 : INV_X1 port map( A => A(14), ZN => n127);
   U135 : OAI21_X1 port map( B1 => SH(4), B2 => n41, A => n3, ZN => B_13_port);
   U136 : AOI221_X1 port map( B1 => n74, B2 => n73, C1 => n70, C2 => n75, A => 
                           n141, ZN => n41);
   U137 : INV_X1 port map( A => n142, ZN => n141);
   U138 : AOI22_X1 port map( A1 => n136, A2 => n79, B1 => n78, B2 => n72, ZN =>
                           n142);
   U139 : OAI221_X1 port map( B1 => n33, B2 => n143, C1 => n34, C2 => n144, A 
                           => n145, ZN => n72);
   U140 : AOI22_X1 port map( A1 => A(3), A2 => n37, B1 => A(2), B2 => n38, ZN 
                           => n145);
   U141 : INV_X1 port map( A => A(4), ZN => n143);
   U142 : MUX2_X1 port map( A => A(1), B => A(0), S => n34, Z => n79);
   U143 : AND2_X1 port map( A1 => SH(2), A2 => SH(3), ZN => n136);
   U144 : OAI221_X1 port map( B1 => n33, B2 => n146, C1 => n34, C2 => n133, A 
                           => n147, ZN => n70);
   U145 : AOI22_X1 port map( A1 => A(11), A2 => n37, B1 => A(10), B2 => n38, ZN
                           => n147);
   U146 : INV_X1 port map( A => A(13), ZN => n133);
   U147 : OAI221_X1 port map( B1 => n33, B2 => n148, C1 => n34, C2 => n149, A 
                           => n150, ZN => n74);
   U148 : AOI22_X1 port map( A1 => A(7), A2 => n37, B1 => A(6), B2 => n38, ZN 
                           => n150);
   U149 : OAI21_X1 port map( B1 => SH(4), B2 => n48, A => n3, ZN => B_12_port);
   U150 : AOI221_X1 port map( B1 => n87, B2 => n73, C1 => n84, C2 => n75, A => 
                           n151, ZN => n48);
   U151 : INV_X1 port map( A => n152, ZN => n151);
   U152 : AOI21_X1 port map( B1 => n78, B2 => n86, A => n80, ZN => n152);
   U153 : OAI221_X1 port map( B1 => n20, B2 => n153, C1 => n154, C2 => n22, A 
                           => n155, ZN => n86);
   U154 : AOI22_X1 port map( A1 => n25, A2 => A(3), B1 => A(4), B2 => n26, ZN 
                           => n155);
   U155 : OAI221_X1 port map( B1 => n33, B2 => n156, C1 => n34, C2 => n146, A 
                           => n157, ZN => n84);
   U156 : AOI22_X1 port map( A1 => A(10), A2 => n37, B1 => A(9), B2 => n38, ZN 
                           => n157);
   U157 : INV_X1 port map( A => A(12), ZN => n146);
   U158 : OAI221_X1 port map( B1 => n33, B2 => n158, C1 => n34, C2 => n148, A 
                           => n159, ZN => n87);
   U159 : AOI22_X1 port map( A1 => A(6), A2 => n37, B1 => A(5), B2 => n38, ZN 
                           => n159);
   U160 : INV_X1 port map( A => A(8), ZN => n148);
   U161 : OAI21_X1 port map( B1 => SH(4), B2 => n56, A => n3, ZN => B_11_port);
   U162 : AOI221_X1 port map( B1 => n95, B2 => n73, C1 => n92, C2 => n75, A => 
                           n160, ZN => n56);
   U163 : INV_X1 port map( A => n161, ZN => n160);
   U164 : AOI21_X1 port map( B1 => n78, B2 => n94, A => n80, ZN => n161);
   U165 : OAI221_X1 port map( B1 => n154, B2 => n20, C1 => n124, C2 => n22, A 
                           => n162, ZN => n94);
   U166 : AOI22_X1 port map( A1 => n25, A2 => A(2), B1 => A(3), B2 => n26, ZN 
                           => n162);
   U167 : INV_X1 port map( A => n34, ZN => n26);
   U168 : INV_X1 port map( A => n33, ZN => n25);
   U169 : OAI221_X1 port map( B1 => n33, B2 => n163, C1 => n34, C2 => n156, A 
                           => n164, ZN => n92);
   U170 : AOI22_X1 port map( A1 => A(9), A2 => n37, B1 => A(8), B2 => n38, ZN 
                           => n164);
   U171 : INV_X1 port map( A => A(11), ZN => n156);
   U172 : OAI221_X1 port map( B1 => n33, B2 => n165, C1 => n34, C2 => n158, A 
                           => n166, ZN => n95);
   U173 : AOI22_X1 port map( A1 => A(5), A2 => n37, B1 => A(4), B2 => n38, ZN 
                           => n166);
   U174 : INV_X1 port map( A => A(7), ZN => n158);
   U175 : OAI21_X1 port map( B1 => SH(4), B2 => n63, A => n3, ZN => B_10_port);
   U176 : NAND2_X1 port map( A1 => SH(4), A2 => A(0), ZN => n3);
   U177 : AOI221_X1 port map( B1 => n102, B2 => n73, C1 => n99, C2 => n75, A =>
                           n167, ZN => n63);
   U178 : INV_X1 port map( A => n168, ZN => n167);
   U179 : AOI21_X1 port map( B1 => n78, B2 => n101, A => n80, ZN => n168);
   U180 : NOR2_X1 port map( A1 => n125, A2 => n107, ZN => n80);
   U181 : NAND2_X1 port map( A1 => SH(3), A2 => A(0), ZN => n107);
   U182 : OAI222_X1 port map( A1 => n34, A2 => n153, B1 => n154, B2 => n33, C1 
                           => n124, C2 => n169, ZN => n101);
   U183 : INV_X1 port map( A => A(0), ZN => n124);
   U184 : INV_X1 port map( A => A(1), ZN => n154);
   U185 : INV_X1 port map( A => A(2), ZN => n153);
   U186 : AND2_X1 port map( A1 => SH(3), A2 => n125, ZN => n78);
   U187 : OAI221_X1 port map( B1 => n33, B2 => n149, C1 => n34, C2 => n163, A 
                           => n170, ZN => n99);
   U188 : AOI22_X1 port map( A1 => A(8), A2 => n37, B1 => A(7), B2 => n38, ZN 
                           => n170);
   U189 : INV_X1 port map( A => A(10), ZN => n163);
   U190 : INV_X1 port map( A => A(9), ZN => n149);
   U191 : NOR2_X1 port map( A1 => n125, A2 => SH(3), ZN => n73);
   U192 : INV_X1 port map( A => SH(2), ZN => n125);
   U193 : INV_X1 port map( A => n171, ZN => n102);
   U194 : AOI221_X1 port map( B1 => n37, B2 => A(4), C1 => A(3), C2 => n38, A 
                           => n172, ZN => n171);
   U195 : OAI22_X1 port map( A1 => n144, A2 => n33, B1 => n165, B2 => n34, ZN 
                           => n172);
   U196 : NAND2_X1 port map( A1 => n173, A2 => n169, ZN => n34);
   U197 : INV_X1 port map( A => A(6), ZN => n165);
   U198 : NAND2_X1 port map( A1 => SH(0), A2 => n169, ZN => n33);
   U199 : INV_X1 port map( A => SH(1), ZN => n169);
   U200 : INV_X1 port map( A => A(5), ZN => n144);
   U201 : INV_X1 port map( A => n22, ZN => n38);
   U202 : NAND2_X1 port map( A1 => SH(0), A2 => SH(1), ZN => n22);
   U203 : INV_X1 port map( A => n20, ZN => n37);
   U204 : NAND2_X1 port map( A1 => SH(1), A2 => n173, ZN => n20);
   U205 : INV_X1 port map( A => SH(0), ZN => n173);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32_DW01_ash_0 is

   port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH : 
         in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out 
         std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32_DW01_ash_0;

architecture SYN_mx2 of SHIFTER_GENERIC_N32_DW01_ash_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   signal SHMAG_3_port, SHMAG_2_port, SHMAG_1_port, SHMAG_0_port, 
      ML_int_1_31_port, ML_int_1_30_port, ML_int_1_29_port, ML_int_1_28_port, 
      ML_int_1_27_port, ML_int_1_26_port, ML_int_1_25_port, ML_int_1_24_port, 
      ML_int_1_23_port, ML_int_1_22_port, ML_int_1_21_port, ML_int_1_20_port, 
      ML_int_1_19_port, ML_int_1_18_port, ML_int_1_17_port, ML_int_1_16_port, 
      ML_int_1_15_port, ML_int_1_14_port, ML_int_1_13_port, ML_int_1_12_port, 
      ML_int_1_11_port, ML_int_1_10_port, ML_int_1_9_port, ML_int_1_8_port, 
      ML_int_1_7_port, ML_int_1_6_port, ML_int_1_5_port, ML_int_1_4_port, 
      ML_int_1_3_port, ML_int_1_2_port, ML_int_1_1_port, ML_int_1_0_port, 
      ML_int_2_31_port, ML_int_2_30_port, ML_int_2_29_port, ML_int_2_28_port, 
      ML_int_2_27_port, ML_int_2_26_port, ML_int_2_25_port, ML_int_2_24_port, 
      ML_int_2_23_port, ML_int_2_22_port, ML_int_2_21_port, ML_int_2_20_port, 
      ML_int_2_19_port, ML_int_2_18_port, ML_int_2_17_port, ML_int_2_16_port, 
      ML_int_2_15_port, ML_int_2_14_port, ML_int_2_13_port, ML_int_2_12_port, 
      ML_int_2_11_port, ML_int_2_10_port, ML_int_2_9_port, ML_int_2_8_port, 
      ML_int_2_7_port, ML_int_2_6_port, ML_int_2_5_port, ML_int_2_4_port, 
      ML_int_2_3_port, ML_int_2_2_port, ML_int_2_1_port, ML_int_2_0_port, 
      ML_int_3_31_port, ML_int_3_30_port, ML_int_3_29_port, ML_int_3_28_port, 
      ML_int_3_27_port, ML_int_3_26_port, ML_int_3_25_port, ML_int_3_24_port, 
      ML_int_3_23_port, ML_int_3_22_port, ML_int_3_21_port, ML_int_3_20_port, 
      ML_int_3_19_port, ML_int_3_18_port, ML_int_3_17_port, ML_int_3_16_port, 
      ML_int_3_15_port, ML_int_3_14_port, ML_int_3_13_port, ML_int_3_12_port, 
      ML_int_3_11_port, ML_int_3_10_port, ML_int_3_9_port, ML_int_3_8_port, 
      ML_int_3_7_port, ML_int_3_6_port, ML_int_3_5_port, ML_int_3_4_port, 
      ML_int_3_3_port, ML_int_3_2_port, ML_int_3_1_port, ML_int_3_0_port, 
      ML_int_4_31_port, ML_int_4_30_port, ML_int_4_29_port, ML_int_4_28_port, 
      ML_int_4_27_port, ML_int_4_26_port, ML_int_4_25_port, ML_int_4_24_port, 
      ML_int_4_23_port, ML_int_4_22_port, ML_int_4_21_port, ML_int_4_20_port, 
      ML_int_4_19_port, ML_int_4_18_port, ML_int_4_17_port, ML_int_4_16_port, 
      ML_int_4_15_port, ML_int_4_14_port, ML_int_4_13_port, ML_int_4_12_port, 
      ML_int_4_11_port, ML_int_4_10_port, ML_int_4_9_port, ML_int_4_8_port, 
      ML_int_4_7_port, ML_int_4_6_port, ML_int_4_5_port, ML_int_4_4_port, 
      ML_int_4_3_port, ML_int_4_2_port, ML_int_4_1_port, ML_int_4_0_port, n1, 
      n2, n3, n4, n5, n6, n7, n8, n9, n10 : std_logic;

begin
   
   M1_4_31 : MUX2_X1 port map( A => ML_int_4_31_port, B => ML_int_4_15_port, S 
                           => n1, Z => B(31));
   M1_4_30 : MUX2_X1 port map( A => ML_int_4_30_port, B => ML_int_4_14_port, S 
                           => n1, Z => B(30));
   M1_4_29 : MUX2_X1 port map( A => ML_int_4_29_port, B => ML_int_4_13_port, S 
                           => n1, Z => B(29));
   M1_4_28 : MUX2_X1 port map( A => ML_int_4_28_port, B => ML_int_4_12_port, S 
                           => n1, Z => B(28));
   M1_4_27 : MUX2_X1 port map( A => ML_int_4_27_port, B => ML_int_4_11_port, S 
                           => n1, Z => B(27));
   M1_4_26 : MUX2_X1 port map( A => ML_int_4_26_port, B => ML_int_4_10_port, S 
                           => n1, Z => B(26));
   M1_4_25 : MUX2_X1 port map( A => ML_int_4_25_port, B => ML_int_4_9_port, S 
                           => n1, Z => B(25));
   M1_4_24 : MUX2_X1 port map( A => ML_int_4_24_port, B => ML_int_4_8_port, S 
                           => n1, Z => B(24));
   M1_4_23 : MUX2_X1 port map( A => ML_int_4_23_port, B => ML_int_4_7_port, S 
                           => n1, Z => B(23));
   M1_4_22 : MUX2_X1 port map( A => ML_int_4_22_port, B => ML_int_4_6_port, S 
                           => n1, Z => B(22));
   M1_4_21 : MUX2_X1 port map( A => ML_int_4_21_port, B => ML_int_4_5_port, S 
                           => n1, Z => B(21));
   M1_4_20 : MUX2_X1 port map( A => ML_int_4_20_port, B => ML_int_4_4_port, S 
                           => n1, Z => B(20));
   M1_4_19 : MUX2_X1 port map( A => ML_int_4_19_port, B => ML_int_4_3_port, S 
                           => n1, Z => B(19));
   M1_4_18 : MUX2_X1 port map( A => ML_int_4_18_port, B => ML_int_4_2_port, S 
                           => n1, Z => B(18));
   M1_4_17 : MUX2_X1 port map( A => ML_int_4_17_port, B => ML_int_4_1_port, S 
                           => n1, Z => B(17));
   M1_4_16 : MUX2_X1 port map( A => ML_int_4_16_port, B => ML_int_4_0_port, S 
                           => n1, Z => B(16));
   M1_3_31 : MUX2_X1 port map( A => ML_int_3_31_port, B => ML_int_3_23_port, S 
                           => SH(3), Z => ML_int_4_31_port);
   M1_3_30 : MUX2_X1 port map( A => ML_int_3_30_port, B => ML_int_3_22_port, S 
                           => SH(3), Z => ML_int_4_30_port);
   M1_3_29 : MUX2_X1 port map( A => ML_int_3_29_port, B => ML_int_3_21_port, S 
                           => SH(3), Z => ML_int_4_29_port);
   M1_3_28 : MUX2_X1 port map( A => ML_int_3_28_port, B => ML_int_3_20_port, S 
                           => SH(3), Z => ML_int_4_28_port);
   M1_3_27 : MUX2_X1 port map( A => ML_int_3_27_port, B => ML_int_3_19_port, S 
                           => SH(3), Z => ML_int_4_27_port);
   M1_3_26 : MUX2_X1 port map( A => ML_int_3_26_port, B => ML_int_3_18_port, S 
                           => SH(3), Z => ML_int_4_26_port);
   M1_3_25 : MUX2_X1 port map( A => ML_int_3_25_port, B => ML_int_3_17_port, S 
                           => SH(3), Z => ML_int_4_25_port);
   M1_3_24 : MUX2_X1 port map( A => ML_int_3_24_port, B => ML_int_3_16_port, S 
                           => SH(3), Z => ML_int_4_24_port);
   M1_3_23 : MUX2_X1 port map( A => ML_int_3_23_port, B => ML_int_3_15_port, S 
                           => SH(3), Z => ML_int_4_23_port);
   M1_3_22 : MUX2_X1 port map( A => ML_int_3_22_port, B => ML_int_3_14_port, S 
                           => SH(3), Z => ML_int_4_22_port);
   M1_3_21 : MUX2_X1 port map( A => ML_int_3_21_port, B => ML_int_3_13_port, S 
                           => SH(3), Z => ML_int_4_21_port);
   M1_3_20 : MUX2_X1 port map( A => ML_int_3_20_port, B => ML_int_3_12_port, S 
                           => SH(3), Z => ML_int_4_20_port);
   M1_3_19 : MUX2_X1 port map( A => ML_int_3_19_port, B => ML_int_3_11_port, S 
                           => SH(3), Z => ML_int_4_19_port);
   M1_3_18 : MUX2_X1 port map( A => ML_int_3_18_port, B => ML_int_3_10_port, S 
                           => SH(3), Z => ML_int_4_18_port);
   M1_3_17 : MUX2_X1 port map( A => ML_int_3_17_port, B => ML_int_3_9_port, S 
                           => SH(3), Z => ML_int_4_17_port);
   M1_3_16 : MUX2_X1 port map( A => ML_int_3_16_port, B => ML_int_3_8_port, S 
                           => SH(3), Z => ML_int_4_16_port);
   M1_3_15 : MUX2_X1 port map( A => ML_int_3_15_port, B => ML_int_3_7_port, S 
                           => SH(3), Z => ML_int_4_15_port);
   M1_3_14 : MUX2_X1 port map( A => ML_int_3_14_port, B => ML_int_3_6_port, S 
                           => SH(3), Z => ML_int_4_14_port);
   M1_3_13 : MUX2_X1 port map( A => ML_int_3_13_port, B => ML_int_3_5_port, S 
                           => SH(3), Z => ML_int_4_13_port);
   M1_3_12 : MUX2_X1 port map( A => ML_int_3_12_port, B => ML_int_3_4_port, S 
                           => SH(3), Z => ML_int_4_12_port);
   M1_3_11 : MUX2_X1 port map( A => ML_int_3_11_port, B => ML_int_3_3_port, S 
                           => SH(3), Z => ML_int_4_11_port);
   M1_3_10 : MUX2_X1 port map( A => ML_int_3_10_port, B => ML_int_3_2_port, S 
                           => SH(3), Z => ML_int_4_10_port);
   M1_3_9 : MUX2_X1 port map( A => ML_int_3_9_port, B => ML_int_3_1_port, S => 
                           SH(3), Z => ML_int_4_9_port);
   M1_3_8 : MUX2_X1 port map( A => ML_int_3_8_port, B => ML_int_3_0_port, S => 
                           SH(3), Z => ML_int_4_8_port);
   M1_2_31 : MUX2_X1 port map( A => ML_int_2_31_port, B => ML_int_2_27_port, S 
                           => SH(2), Z => ML_int_3_31_port);
   M1_2_30 : MUX2_X1 port map( A => ML_int_2_30_port, B => ML_int_2_26_port, S 
                           => SH(2), Z => ML_int_3_30_port);
   M1_2_29 : MUX2_X1 port map( A => ML_int_2_29_port, B => ML_int_2_25_port, S 
                           => SH(2), Z => ML_int_3_29_port);
   M1_2_28 : MUX2_X1 port map( A => ML_int_2_28_port, B => ML_int_2_24_port, S 
                           => SH(2), Z => ML_int_3_28_port);
   M1_2_27 : MUX2_X1 port map( A => ML_int_2_27_port, B => ML_int_2_23_port, S 
                           => SH(2), Z => ML_int_3_27_port);
   M1_2_26 : MUX2_X1 port map( A => ML_int_2_26_port, B => ML_int_2_22_port, S 
                           => SH(2), Z => ML_int_3_26_port);
   M1_2_25 : MUX2_X1 port map( A => ML_int_2_25_port, B => ML_int_2_21_port, S 
                           => SH(2), Z => ML_int_3_25_port);
   M1_2_24 : MUX2_X1 port map( A => ML_int_2_24_port, B => ML_int_2_20_port, S 
                           => SH(2), Z => ML_int_3_24_port);
   M1_2_23 : MUX2_X1 port map( A => ML_int_2_23_port, B => ML_int_2_19_port, S 
                           => SH(2), Z => ML_int_3_23_port);
   M1_2_22 : MUX2_X1 port map( A => ML_int_2_22_port, B => ML_int_2_18_port, S 
                           => SH(2), Z => ML_int_3_22_port);
   M1_2_21 : MUX2_X1 port map( A => ML_int_2_21_port, B => ML_int_2_17_port, S 
                           => SH(2), Z => ML_int_3_21_port);
   M1_2_20 : MUX2_X1 port map( A => ML_int_2_20_port, B => ML_int_2_16_port, S 
                           => SH(2), Z => ML_int_3_20_port);
   M1_2_19 : MUX2_X1 port map( A => ML_int_2_19_port, B => ML_int_2_15_port, S 
                           => SH(2), Z => ML_int_3_19_port);
   M1_2_18 : MUX2_X1 port map( A => ML_int_2_18_port, B => ML_int_2_14_port, S 
                           => SH(2), Z => ML_int_3_18_port);
   M1_2_17 : MUX2_X1 port map( A => ML_int_2_17_port, B => ML_int_2_13_port, S 
                           => SH(2), Z => ML_int_3_17_port);
   M1_2_16 : MUX2_X1 port map( A => ML_int_2_16_port, B => ML_int_2_12_port, S 
                           => SH(2), Z => ML_int_3_16_port);
   M1_2_15 : MUX2_X1 port map( A => ML_int_2_15_port, B => ML_int_2_11_port, S 
                           => SH(2), Z => ML_int_3_15_port);
   M1_2_14 : MUX2_X1 port map( A => ML_int_2_14_port, B => ML_int_2_10_port, S 
                           => SH(2), Z => ML_int_3_14_port);
   M1_2_13 : MUX2_X1 port map( A => ML_int_2_13_port, B => ML_int_2_9_port, S 
                           => SH(2), Z => ML_int_3_13_port);
   M1_2_12 : MUX2_X1 port map( A => ML_int_2_12_port, B => ML_int_2_8_port, S 
                           => SH(2), Z => ML_int_3_12_port);
   M1_2_11 : MUX2_X1 port map( A => ML_int_2_11_port, B => ML_int_2_7_port, S 
                           => SH(2), Z => ML_int_3_11_port);
   M1_2_10 : MUX2_X1 port map( A => ML_int_2_10_port, B => ML_int_2_6_port, S 
                           => SH(2), Z => ML_int_3_10_port);
   M1_2_9 : MUX2_X1 port map( A => ML_int_2_9_port, B => ML_int_2_5_port, S => 
                           SH(2), Z => ML_int_3_9_port);
   M1_2_8 : MUX2_X1 port map( A => ML_int_2_8_port, B => ML_int_2_4_port, S => 
                           SH(2), Z => ML_int_3_8_port);
   M1_2_7 : MUX2_X1 port map( A => ML_int_2_7_port, B => ML_int_2_3_port, S => 
                           SH(2), Z => ML_int_3_7_port);
   M1_2_6 : MUX2_X1 port map( A => ML_int_2_6_port, B => ML_int_2_2_port, S => 
                           SH(2), Z => ML_int_3_6_port);
   M1_2_5 : MUX2_X1 port map( A => ML_int_2_5_port, B => ML_int_2_1_port, S => 
                           SH(2), Z => ML_int_3_5_port);
   M1_2_4 : MUX2_X1 port map( A => ML_int_2_4_port, B => ML_int_2_0_port, S => 
                           SH(2), Z => ML_int_3_4_port);
   M1_1_31 : MUX2_X1 port map( A => ML_int_1_31_port, B => ML_int_1_29_port, S 
                           => SH(1), Z => ML_int_2_31_port);
   M1_1_30 : MUX2_X1 port map( A => ML_int_1_30_port, B => ML_int_1_28_port, S 
                           => SH(1), Z => ML_int_2_30_port);
   M1_1_29 : MUX2_X1 port map( A => ML_int_1_29_port, B => ML_int_1_27_port, S 
                           => SH(1), Z => ML_int_2_29_port);
   M1_1_28 : MUX2_X1 port map( A => ML_int_1_28_port, B => ML_int_1_26_port, S 
                           => SH(1), Z => ML_int_2_28_port);
   M1_1_27 : MUX2_X1 port map( A => ML_int_1_27_port, B => ML_int_1_25_port, S 
                           => SH(1), Z => ML_int_2_27_port);
   M1_1_26 : MUX2_X1 port map( A => ML_int_1_26_port, B => ML_int_1_24_port, S 
                           => SH(1), Z => ML_int_2_26_port);
   M1_1_25 : MUX2_X1 port map( A => ML_int_1_25_port, B => ML_int_1_23_port, S 
                           => SH(1), Z => ML_int_2_25_port);
   M1_1_24 : MUX2_X1 port map( A => ML_int_1_24_port, B => ML_int_1_22_port, S 
                           => SH(1), Z => ML_int_2_24_port);
   M1_1_23 : MUX2_X1 port map( A => ML_int_1_23_port, B => ML_int_1_21_port, S 
                           => SH(1), Z => ML_int_2_23_port);
   M1_1_22 : MUX2_X1 port map( A => ML_int_1_22_port, B => ML_int_1_20_port, S 
                           => SH(1), Z => ML_int_2_22_port);
   M1_1_21 : MUX2_X1 port map( A => ML_int_1_21_port, B => ML_int_1_19_port, S 
                           => SH(1), Z => ML_int_2_21_port);
   M1_1_20 : MUX2_X1 port map( A => ML_int_1_20_port, B => ML_int_1_18_port, S 
                           => SH(1), Z => ML_int_2_20_port);
   M1_1_19 : MUX2_X1 port map( A => ML_int_1_19_port, B => ML_int_1_17_port, S 
                           => SH(1), Z => ML_int_2_19_port);
   M1_1_18 : MUX2_X1 port map( A => ML_int_1_18_port, B => ML_int_1_16_port, S 
                           => SH(1), Z => ML_int_2_18_port);
   M1_1_17 : MUX2_X1 port map( A => ML_int_1_17_port, B => ML_int_1_15_port, S 
                           => SH(1), Z => ML_int_2_17_port);
   M1_1_16 : MUX2_X1 port map( A => ML_int_1_16_port, B => ML_int_1_14_port, S 
                           => SH(1), Z => ML_int_2_16_port);
   M1_1_15 : MUX2_X1 port map( A => ML_int_1_15_port, B => ML_int_1_13_port, S 
                           => SH(1), Z => ML_int_2_15_port);
   M1_1_14 : MUX2_X1 port map( A => ML_int_1_14_port, B => ML_int_1_12_port, S 
                           => SH(1), Z => ML_int_2_14_port);
   M1_1_13 : MUX2_X1 port map( A => ML_int_1_13_port, B => ML_int_1_11_port, S 
                           => SH(1), Z => ML_int_2_13_port);
   M1_1_12 : MUX2_X1 port map( A => ML_int_1_12_port, B => ML_int_1_10_port, S 
                           => SH(1), Z => ML_int_2_12_port);
   M1_1_11 : MUX2_X1 port map( A => ML_int_1_11_port, B => ML_int_1_9_port, S 
                           => SH(1), Z => ML_int_2_11_port);
   M1_1_10 : MUX2_X1 port map( A => ML_int_1_10_port, B => ML_int_1_8_port, S 
                           => SH(1), Z => ML_int_2_10_port);
   M1_1_9 : MUX2_X1 port map( A => ML_int_1_9_port, B => ML_int_1_7_port, S => 
                           SH(1), Z => ML_int_2_9_port);
   M1_1_8 : MUX2_X1 port map( A => ML_int_1_8_port, B => ML_int_1_6_port, S => 
                           SH(1), Z => ML_int_2_8_port);
   M1_1_7 : MUX2_X1 port map( A => ML_int_1_7_port, B => ML_int_1_5_port, S => 
                           SH(1), Z => ML_int_2_7_port);
   M1_1_6 : MUX2_X1 port map( A => ML_int_1_6_port, B => ML_int_1_4_port, S => 
                           SH(1), Z => ML_int_2_6_port);
   M1_1_5 : MUX2_X1 port map( A => ML_int_1_5_port, B => ML_int_1_3_port, S => 
                           SH(1), Z => ML_int_2_5_port);
   M1_1_4 : MUX2_X1 port map( A => ML_int_1_4_port, B => ML_int_1_2_port, S => 
                           SH(1), Z => ML_int_2_4_port);
   M1_1_3 : MUX2_X1 port map( A => ML_int_1_3_port, B => ML_int_1_1_port, S => 
                           SH(1), Z => ML_int_2_3_port);
   M1_1_2 : MUX2_X1 port map( A => ML_int_1_2_port, B => ML_int_1_0_port, S => 
                           SH(1), Z => ML_int_2_2_port);
   M1_0_31 : MUX2_X1 port map( A => A(31), B => A(30), S => SH(0), Z => 
                           ML_int_1_31_port);
   M1_0_30 : MUX2_X1 port map( A => A(30), B => A(29), S => SH(0), Z => 
                           ML_int_1_30_port);
   M1_0_29 : MUX2_X1 port map( A => A(29), B => A(28), S => SH(0), Z => 
                           ML_int_1_29_port);
   M1_0_28 : MUX2_X1 port map( A => A(28), B => A(27), S => SH(0), Z => 
                           ML_int_1_28_port);
   M1_0_27 : MUX2_X1 port map( A => A(27), B => A(26), S => SH(0), Z => 
                           ML_int_1_27_port);
   M1_0_26 : MUX2_X1 port map( A => A(26), B => A(25), S => SH(0), Z => 
                           ML_int_1_26_port);
   M1_0_25 : MUX2_X1 port map( A => A(25), B => A(24), S => SH(0), Z => 
                           ML_int_1_25_port);
   M1_0_24 : MUX2_X1 port map( A => A(24), B => A(23), S => SH(0), Z => 
                           ML_int_1_24_port);
   M1_0_23 : MUX2_X1 port map( A => A(23), B => A(22), S => SH(0), Z => 
                           ML_int_1_23_port);
   M1_0_22 : MUX2_X1 port map( A => A(22), B => A(21), S => SH(0), Z => 
                           ML_int_1_22_port);
   M1_0_21 : MUX2_X1 port map( A => A(21), B => A(20), S => SH(0), Z => 
                           ML_int_1_21_port);
   M1_0_20 : MUX2_X1 port map( A => A(20), B => A(19), S => SH(0), Z => 
                           ML_int_1_20_port);
   M1_0_19 : MUX2_X1 port map( A => A(19), B => A(18), S => SH(0), Z => 
                           ML_int_1_19_port);
   M1_0_18 : MUX2_X1 port map( A => A(18), B => A(17), S => SH(0), Z => 
                           ML_int_1_18_port);
   M1_0_17 : MUX2_X1 port map( A => A(17), B => A(16), S => SH(0), Z => 
                           ML_int_1_17_port);
   M1_0_16 : MUX2_X1 port map( A => A(16), B => A(15), S => SH(0), Z => 
                           ML_int_1_16_port);
   M1_0_15 : MUX2_X1 port map( A => A(15), B => A(14), S => SH(0), Z => 
                           ML_int_1_15_port);
   M1_0_14 : MUX2_X1 port map( A => A(14), B => A(13), S => SH(0), Z => 
                           ML_int_1_14_port);
   M1_0_13 : MUX2_X1 port map( A => A(13), B => A(12), S => SH(0), Z => 
                           ML_int_1_13_port);
   M1_0_12 : MUX2_X1 port map( A => A(12), B => A(11), S => SH(0), Z => 
                           ML_int_1_12_port);
   M1_0_11 : MUX2_X1 port map( A => A(11), B => A(10), S => SH(0), Z => 
                           ML_int_1_11_port);
   M1_0_10 : MUX2_X1 port map( A => A(10), B => A(9), S => SH(0), Z => 
                           ML_int_1_10_port);
   M1_0_9 : MUX2_X1 port map( A => A(9), B => A(8), S => SH(0), Z => 
                           ML_int_1_9_port);
   M1_0_8 : MUX2_X1 port map( A => A(8), B => A(7), S => SH(0), Z => 
                           ML_int_1_8_port);
   M1_0_7 : MUX2_X1 port map( A => A(7), B => A(6), S => SH(0), Z => 
                           ML_int_1_7_port);
   M1_0_6 : MUX2_X1 port map( A => A(6), B => A(5), S => SH(0), Z => 
                           ML_int_1_6_port);
   M1_0_5 : MUX2_X1 port map( A => A(5), B => A(4), S => SH(0), Z => 
                           ML_int_1_5_port);
   M1_0_4 : MUX2_X1 port map( A => A(4), B => A(3), S => SH(0), Z => 
                           ML_int_1_4_port);
   M1_0_3 : MUX2_X1 port map( A => A(3), B => A(2), S => SH(0), Z => 
                           ML_int_1_3_port);
   M1_0_2 : MUX2_X1 port map( A => A(2), B => A(1), S => SH(0), Z => 
                           ML_int_1_2_port);
   M1_0_1 : MUX2_X1 port map( A => A(1), B => A(0), S => SH(0), Z => 
                           ML_int_1_1_port);
   U3 : INV_X1 port map( A => n2, ZN => n1);
   U4 : INV_X1 port map( A => SH(4), ZN => n2);
   U5 : AND2_X1 port map( A1 => ML_int_4_9_port, A2 => n2, ZN => B(9));
   U6 : AND2_X1 port map( A1 => ML_int_4_8_port, A2 => n2, ZN => B(8));
   U7 : NOR2_X1 port map( A1 => n1, A2 => n3, ZN => B(7));
   U8 : NOR2_X1 port map( A1 => n1, A2 => n4, ZN => B(6));
   U9 : NOR2_X1 port map( A1 => n1, A2 => n5, ZN => B(5));
   U10 : NOR2_X1 port map( A1 => n1, A2 => n6, ZN => B(4));
   U11 : NOR2_X1 port map( A1 => n1, A2 => n7, ZN => B(3));
   U12 : NOR2_X1 port map( A1 => n1, A2 => n8, ZN => B(2));
   U13 : NOR2_X1 port map( A1 => n1, A2 => n9, ZN => B(1));
   U14 : AND2_X1 port map( A1 => ML_int_4_15_port, A2 => n2, ZN => B(15));
   U15 : AND2_X1 port map( A1 => ML_int_4_14_port, A2 => n2, ZN => B(14));
   U16 : AND2_X1 port map( A1 => ML_int_4_13_port, A2 => n2, ZN => B(13));
   U17 : AND2_X1 port map( A1 => ML_int_4_12_port, A2 => n2, ZN => B(12));
   U18 : AND2_X1 port map( A1 => ML_int_4_11_port, A2 => n2, ZN => B(11));
   U19 : AND2_X1 port map( A1 => ML_int_4_10_port, A2 => n2, ZN => B(10));
   U20 : NOR2_X1 port map( A1 => SH(4), A2 => n10, ZN => B(0));
   U21 : INV_X1 port map( A => n3, ZN => ML_int_4_7_port);
   U22 : NAND2_X1 port map( A1 => ML_int_3_7_port, A2 => SHMAG_3_port, ZN => n3
                           );
   U23 : INV_X1 port map( A => n4, ZN => ML_int_4_6_port);
   U24 : NAND2_X1 port map( A1 => ML_int_3_6_port, A2 => SHMAG_3_port, ZN => n4
                           );
   U25 : INV_X1 port map( A => n5, ZN => ML_int_4_5_port);
   U26 : NAND2_X1 port map( A1 => ML_int_3_5_port, A2 => SHMAG_3_port, ZN => n5
                           );
   U27 : INV_X1 port map( A => n6, ZN => ML_int_4_4_port);
   U28 : NAND2_X1 port map( A1 => ML_int_3_4_port, A2 => SHMAG_3_port, ZN => n6
                           );
   U29 : INV_X1 port map( A => n7, ZN => ML_int_4_3_port);
   U30 : NAND2_X1 port map( A1 => ML_int_3_3_port, A2 => SHMAG_3_port, ZN => n7
                           );
   U31 : INV_X1 port map( A => n8, ZN => ML_int_4_2_port);
   U32 : NAND2_X1 port map( A1 => ML_int_3_2_port, A2 => SHMAG_3_port, ZN => n8
                           );
   U33 : INV_X1 port map( A => n9, ZN => ML_int_4_1_port);
   U34 : NAND2_X1 port map( A1 => ML_int_3_1_port, A2 => SHMAG_3_port, ZN => n9
                           );
   U35 : INV_X1 port map( A => n10, ZN => ML_int_4_0_port);
   U36 : NAND2_X1 port map( A1 => ML_int_3_0_port, A2 => SHMAG_3_port, ZN => 
                           n10);
   U37 : INV_X1 port map( A => SH(3), ZN => SHMAG_3_port);
   U38 : AND2_X1 port map( A1 => ML_int_2_3_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_3_port);
   U39 : AND2_X1 port map( A1 => ML_int_2_2_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_2_port);
   U40 : AND2_X1 port map( A1 => ML_int_2_1_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_1_port);
   U41 : AND2_X1 port map( A1 => ML_int_2_0_port, A2 => SHMAG_2_port, ZN => 
                           ML_int_3_0_port);
   U42 : INV_X1 port map( A => SH(2), ZN => SHMAG_2_port);
   U43 : AND2_X1 port map( A1 => ML_int_1_1_port, A2 => SHMAG_1_port, ZN => 
                           ML_int_2_1_port);
   U44 : AND2_X1 port map( A1 => ML_int_1_0_port, A2 => SHMAG_1_port, ZN => 
                           ML_int_2_0_port);
   U45 : INV_X1 port map( A => SH(1), ZN => SHMAG_1_port);
   U46 : AND2_X1 port map( A1 => A(0), A2 => SHMAG_0_port, ZN => 
                           ML_int_1_0_port);
   U47 : INV_X1 port map( A => SH(0), ZN => SHMAG_0_port);

end SYN_mx2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32_DW01_add_1 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end DLX_IR_SIZE32_PC_SIZE32_DW01_add_1;

architecture SYN_rpl of DLX_IR_SIZE32_PC_SIZE32_DW01_add_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, carry_31_port, 
      carry_30_port, carry_29_port, carry_28_port, carry_27_port, carry_26_port
      , carry_25_port, carry_24_port, carry_23_port, carry_22_port, 
      carry_21_port, carry_20_port, carry_19_port, carry_18_port, carry_17_port
      , carry_16_port, carry_15_port, carry_14_port, carry_13_port, 
      carry_12_port, carry_11_port, carry_10_port, carry_9_port, carry_8_port, 
      carry_7_port, carry_6_port, carry_5_port, carry_4_port : std_logic;

begin
   SUM <= ( SUM_31_port, SUM_30_port, SUM_29_port, SUM_28_port, SUM_27_port, 
      SUM_26_port, SUM_25_port, SUM_24_port, SUM_23_port, SUM_22_port, 
      SUM_21_port, SUM_20_port, SUM_19_port, SUM_18_port, SUM_17_port, 
      SUM_16_port, SUM_15_port, SUM_14_port, SUM_13_port, SUM_12_port, 
      SUM_11_port, SUM_10_port, SUM_9_port, SUM_8_port, SUM_7_port, SUM_6_port,
      SUM_5_port, SUM_4_port, SUM_3_port, SUM_2_port, A(1), A(0) );
   
   U1 : XOR2_X1 port map( A => A(31), B => carry_31_port, Z => SUM_31_port);
   U2 : AND2_X1 port map( A1 => carry_30_port, A2 => A(30), ZN => carry_31_port
                           );
   U3 : XOR2_X1 port map( A => A(30), B => carry_30_port, Z => SUM_30_port);
   U4 : AND2_X1 port map( A1 => carry_29_port, A2 => A(29), ZN => carry_30_port
                           );
   U5 : XOR2_X1 port map( A => A(29), B => carry_29_port, Z => SUM_29_port);
   U6 : AND2_X1 port map( A1 => carry_28_port, A2 => A(28), ZN => carry_29_port
                           );
   U7 : XOR2_X1 port map( A => A(28), B => carry_28_port, Z => SUM_28_port);
   U8 : AND2_X1 port map( A1 => carry_27_port, A2 => A(27), ZN => carry_28_port
                           );
   U9 : XOR2_X1 port map( A => A(27), B => carry_27_port, Z => SUM_27_port);
   U10 : AND2_X1 port map( A1 => carry_26_port, A2 => A(26), ZN => 
                           carry_27_port);
   U11 : XOR2_X1 port map( A => A(26), B => carry_26_port, Z => SUM_26_port);
   U12 : AND2_X1 port map( A1 => carry_25_port, A2 => A(25), ZN => 
                           carry_26_port);
   U13 : XOR2_X1 port map( A => A(25), B => carry_25_port, Z => SUM_25_port);
   U14 : AND2_X1 port map( A1 => carry_24_port, A2 => A(24), ZN => 
                           carry_25_port);
   U15 : XOR2_X1 port map( A => A(24), B => carry_24_port, Z => SUM_24_port);
   U16 : AND2_X1 port map( A1 => carry_23_port, A2 => A(23), ZN => 
                           carry_24_port);
   U17 : XOR2_X1 port map( A => A(23), B => carry_23_port, Z => SUM_23_port);
   U18 : AND2_X1 port map( A1 => carry_22_port, A2 => A(22), ZN => 
                           carry_23_port);
   U19 : XOR2_X1 port map( A => A(22), B => carry_22_port, Z => SUM_22_port);
   U20 : AND2_X1 port map( A1 => carry_21_port, A2 => A(21), ZN => 
                           carry_22_port);
   U21 : XOR2_X1 port map( A => A(21), B => carry_21_port, Z => SUM_21_port);
   U22 : AND2_X1 port map( A1 => carry_20_port, A2 => A(20), ZN => 
                           carry_21_port);
   U23 : XOR2_X1 port map( A => A(20), B => carry_20_port, Z => SUM_20_port);
   U24 : AND2_X1 port map( A1 => carry_19_port, A2 => A(19), ZN => 
                           carry_20_port);
   U25 : XOR2_X1 port map( A => A(19), B => carry_19_port, Z => SUM_19_port);
   U26 : AND2_X1 port map( A1 => carry_18_port, A2 => A(18), ZN => 
                           carry_19_port);
   U27 : XOR2_X1 port map( A => A(18), B => carry_18_port, Z => SUM_18_port);
   U28 : AND2_X1 port map( A1 => carry_17_port, A2 => A(17), ZN => 
                           carry_18_port);
   U29 : XOR2_X1 port map( A => A(17), B => carry_17_port, Z => SUM_17_port);
   U30 : AND2_X1 port map( A1 => carry_16_port, A2 => A(16), ZN => 
                           carry_17_port);
   U31 : XOR2_X1 port map( A => A(16), B => carry_16_port, Z => SUM_16_port);
   U32 : AND2_X1 port map( A1 => carry_15_port, A2 => A(15), ZN => 
                           carry_16_port);
   U33 : XOR2_X1 port map( A => A(15), B => carry_15_port, Z => SUM_15_port);
   U34 : AND2_X1 port map( A1 => carry_14_port, A2 => A(14), ZN => 
                           carry_15_port);
   U35 : XOR2_X1 port map( A => A(14), B => carry_14_port, Z => SUM_14_port);
   U36 : AND2_X1 port map( A1 => carry_13_port, A2 => A(13), ZN => 
                           carry_14_port);
   U37 : XOR2_X1 port map( A => A(13), B => carry_13_port, Z => SUM_13_port);
   U38 : AND2_X1 port map( A1 => carry_12_port, A2 => A(12), ZN => 
                           carry_13_port);
   U39 : XOR2_X1 port map( A => A(12), B => carry_12_port, Z => SUM_12_port);
   U40 : AND2_X1 port map( A1 => carry_11_port, A2 => A(11), ZN => 
                           carry_12_port);
   U41 : XOR2_X1 port map( A => A(11), B => carry_11_port, Z => SUM_11_port);
   U42 : AND2_X1 port map( A1 => carry_10_port, A2 => A(10), ZN => 
                           carry_11_port);
   U43 : XOR2_X1 port map( A => A(10), B => carry_10_port, Z => SUM_10_port);
   U44 : AND2_X1 port map( A1 => carry_9_port, A2 => A(9), ZN => carry_10_port)
                           ;
   U45 : XOR2_X1 port map( A => A(9), B => carry_9_port, Z => SUM_9_port);
   U46 : AND2_X1 port map( A1 => carry_8_port, A2 => A(8), ZN => carry_9_port);
   U47 : XOR2_X1 port map( A => A(8), B => carry_8_port, Z => SUM_8_port);
   U48 : AND2_X1 port map( A1 => carry_7_port, A2 => A(7), ZN => carry_8_port);
   U49 : XOR2_X1 port map( A => A(7), B => carry_7_port, Z => SUM_7_port);
   U50 : AND2_X1 port map( A1 => carry_6_port, A2 => A(6), ZN => carry_7_port);
   U51 : XOR2_X1 port map( A => A(6), B => carry_6_port, Z => SUM_6_port);
   U52 : AND2_X1 port map( A1 => carry_5_port, A2 => A(5), ZN => carry_6_port);
   U53 : XOR2_X1 port map( A => A(5), B => carry_5_port, Z => SUM_5_port);
   U54 : AND2_X1 port map( A1 => carry_4_port, A2 => A(4), ZN => carry_5_port);
   U55 : XOR2_X1 port map( A => A(4), B => carry_4_port, Z => SUM_4_port);
   U56 : AND2_X1 port map( A1 => A(2), A2 => A(3), ZN => carry_4_port);
   U57 : XOR2_X1 port map( A => A(3), B => A(2), Z => SUM_3_port);
   U58 : INV_X1 port map( A => A(2), ZN => SUM_2_port);

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32_DW01_add_0 is

   port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0);  CO : out std_logic);

end DLX_IR_SIZE32_PC_SIZE32_DW01_add_0;

architecture SYN_rpl of DLX_IR_SIZE32_PC_SIZE32_DW01_add_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component FA_X1
      port( A, B, CI : in std_logic;  CO, S : out std_logic);
   end component;
   
   signal carry_31_port, carry_30_port, carry_29_port, carry_28_port, 
      carry_27_port, carry_26_port, carry_25_port, carry_24_port, carry_23_port
      , carry_22_port, carry_21_port, carry_20_port, carry_19_port, 
      carry_18_port, carry_17_port, carry_16_port, carry_15_port, carry_14_port
      , carry_13_port, carry_12_port, carry_11_port, carry_10_port, 
      carry_9_port, carry_8_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, net43517 : 
      std_logic;

begin
   
   U1_31 : FA_X1 port map( A => A(31), B => B(31), CI => carry_31_port, CO => 
                           net43517, S => SUM(31));
   U1_30 : FA_X1 port map( A => A(30), B => B(30), CI => carry_30_port, CO => 
                           carry_31_port, S => SUM(30));
   U1_29 : FA_X1 port map( A => A(29), B => B(29), CI => carry_29_port, CO => 
                           carry_30_port, S => SUM(29));
   U1_28 : FA_X1 port map( A => A(28), B => B(28), CI => carry_28_port, CO => 
                           carry_29_port, S => SUM(28));
   U1_27 : FA_X1 port map( A => A(27), B => B(27), CI => carry_27_port, CO => 
                           carry_28_port, S => SUM(27));
   U1_26 : FA_X1 port map( A => A(26), B => B(26), CI => carry_26_port, CO => 
                           carry_27_port, S => SUM(26));
   U1_25 : FA_X1 port map( A => A(25), B => B(25), CI => carry_25_port, CO => 
                           carry_26_port, S => SUM(25));
   U1_24 : FA_X1 port map( A => A(24), B => B(24), CI => carry_24_port, CO => 
                           carry_25_port, S => SUM(24));
   U1_23 : FA_X1 port map( A => A(23), B => B(23), CI => carry_23_port, CO => 
                           carry_24_port, S => SUM(23));
   U1_22 : FA_X1 port map( A => A(22), B => B(22), CI => carry_22_port, CO => 
                           carry_23_port, S => SUM(22));
   U1_21 : FA_X1 port map( A => A(21), B => B(21), CI => carry_21_port, CO => 
                           carry_22_port, S => SUM(21));
   U1_20 : FA_X1 port map( A => A(20), B => B(20), CI => carry_20_port, CO => 
                           carry_21_port, S => SUM(20));
   U1_19 : FA_X1 port map( A => A(19), B => B(19), CI => carry_19_port, CO => 
                           carry_20_port, S => SUM(19));
   U1_18 : FA_X1 port map( A => A(18), B => B(18), CI => carry_18_port, CO => 
                           carry_19_port, S => SUM(18));
   U1_17 : FA_X1 port map( A => A(17), B => B(17), CI => carry_17_port, CO => 
                           carry_18_port, S => SUM(17));
   U1_16 : FA_X1 port map( A => A(16), B => B(16), CI => carry_16_port, CO => 
                           carry_17_port, S => SUM(16));
   U1_15 : FA_X1 port map( A => A(15), B => B(15), CI => carry_15_port, CO => 
                           carry_16_port, S => SUM(15));
   U1_14 : FA_X1 port map( A => A(14), B => B(14), CI => carry_14_port, CO => 
                           carry_15_port, S => SUM(14));
   U1_13 : FA_X1 port map( A => A(13), B => B(13), CI => carry_13_port, CO => 
                           carry_14_port, S => SUM(13));
   U1_12 : FA_X1 port map( A => A(12), B => B(12), CI => carry_12_port, CO => 
                           carry_13_port, S => SUM(12));
   U1_11 : FA_X1 port map( A => A(11), B => B(11), CI => carry_11_port, CO => 
                           carry_12_port, S => SUM(11));
   U1_10 : FA_X1 port map( A => A(10), B => B(10), CI => carry_10_port, CO => 
                           carry_11_port, S => SUM(10));
   U1_9 : FA_X1 port map( A => A(9), B => B(9), CI => carry_9_port, CO => 
                           carry_10_port, S => SUM(9));
   U1_8 : FA_X1 port map( A => A(8), B => B(8), CI => carry_8_port, CO => 
                           carry_9_port, S => SUM(8));
   U1_7 : FA_X1 port map( A => A(7), B => B(7), CI => carry_7_port, CO => 
                           carry_8_port, S => SUM(7));
   U1_6 : FA_X1 port map( A => A(6), B => B(6), CI => carry_6_port, CO => 
                           carry_7_port, S => SUM(6));
   U1_5 : FA_X1 port map( A => A(5), B => B(5), CI => carry_5_port, CO => 
                           carry_6_port, S => SUM(5));
   U1_4 : FA_X1 port map( A => A(4), B => B(4), CI => carry_4_port, CO => 
                           carry_5_port, S => SUM(4));
   U1_3 : FA_X1 port map( A => A(3), B => B(3), CI => carry_3_port, CO => 
                           carry_4_port, S => SUM(3));
   U1_2 : FA_X1 port map( A => A(2), B => B(2), CI => carry_2_port, CO => 
                           carry_3_port, S => SUM(2));
   U1_1 : FA_X1 port map( A => A(1), B => B(1), CI => carry_1_port, CO => 
                           carry_2_port, S => SUM(1));
   U1 : AND2_X1 port map( A1 => A(0), A2 => B(0), ZN => carry_1_port);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => SUM(0));

end SYN_rpl;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_generic_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end mux21_generic_NBIT4_7;

architecture SYN_behavioural of mux21_generic_NBIT4_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_generic_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end mux21_generic_NBIT4_6;

architecture SYN_behavioural of mux21_generic_NBIT4_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_generic_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end mux21_generic_NBIT4_5;

architecture SYN_behavioural of mux21_generic_NBIT4_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_generic_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end mux21_generic_NBIT4_4;

architecture SYN_behavioural of mux21_generic_NBIT4_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_generic_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end mux21_generic_NBIT4_3;

architecture SYN_behavioural of mux21_generic_NBIT4_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_generic_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end mux21_generic_NBIT4_2;

architecture SYN_behavioural of mux21_generic_NBIT4_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_generic_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end mux21_generic_NBIT4_1;

architecture SYN_behavioural of mux21_generic_NBIT4_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_15 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_15;

architecture SYN_structural of RCA_GEN_NBIT4_15 is

   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_60 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_59 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_58 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_57 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_14 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_14;

architecture SYN_structural of RCA_GEN_NBIT4_14 is

   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_56 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_55 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_54 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_53 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_13 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_13;

architecture SYN_structural of RCA_GEN_NBIT4_13 is

   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_52 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_51 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_50 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_49 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_12 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_12;

architecture SYN_structural of RCA_GEN_NBIT4_12 is

   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_48 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_47 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_46 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_45 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_11 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_11;

architecture SYN_structural of RCA_GEN_NBIT4_11 is

   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_44 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_43 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_42 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_41 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_10 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_10;

architecture SYN_structural of RCA_GEN_NBIT4_10 is

   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_40 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_39 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_38 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_37 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_9 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_9;

architecture SYN_structural of RCA_GEN_NBIT4_9 is

   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_36 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_35 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_34 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_33 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_8 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_8;

architecture SYN_structural of RCA_GEN_NBIT4_8 is

   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_32 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_31 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_30 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_29 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_7;

architecture SYN_structural of RCA_GEN_NBIT4_7 is

   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_28 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_27 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_26 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_25 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_6;

architecture SYN_structural of RCA_GEN_NBIT4_6 is

   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_24 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_23 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_22 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_21 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_5;

architecture SYN_structural of RCA_GEN_NBIT4_5 is

   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_20 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_19 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_18 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_17 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_4;

architecture SYN_structural of RCA_GEN_NBIT4_4 is

   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_16 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_15 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_14 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_13 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_3;

architecture SYN_structural of RCA_GEN_NBIT4_3 is

   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_12 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_11 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_10 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_9 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_2;

architecture SYN_structural of RCA_GEN_NBIT4_2 is

   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_8 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_7 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_6 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_5 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_1;

architecture SYN_structural of RCA_GEN_NBIT4_1 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_4 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_3 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_2 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_1 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_23 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_23;

architecture SYN_beh of PGnet_23 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_22 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_22;

architecture SYN_beh of PGnet_22 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_21 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_21;

architecture SYN_beh of PGnet_21 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_20 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_20;

architecture SYN_beh of PGnet_20 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_19 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_19;

architecture SYN_beh of PGnet_19 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_18 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_18;

architecture SYN_beh of PGnet_18 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_17 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_17;

architecture SYN_beh of PGnet_17 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_16 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_16;

architecture SYN_beh of PGnet_16 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_15 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_15;

architecture SYN_beh of PGnet_15 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_14 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_14;

architecture SYN_beh of PGnet_14 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_13 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_13;

architecture SYN_beh of PGnet_13 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_12 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_12;

architecture SYN_beh of PGnet_12 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_11 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_11;

architecture SYN_beh of PGnet_11 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_10 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_10;

architecture SYN_beh of PGnet_10 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_9 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_9;

architecture SYN_beh of PGnet_9 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_8 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_8;

architecture SYN_beh of PGnet_8 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_7 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_7;

architecture SYN_beh of PGnet_7 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_6 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_6;

architecture SYN_beh of PGnet_6 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_5 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_5;

architecture SYN_beh of PGnet_5 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_4 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_4;

architecture SYN_beh of PGnet_4 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_3 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_3;

architecture SYN_beh of PGnet_3 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_2 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_2;

architecture SYN_beh of PGnet_2 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_1 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_1;

architecture SYN_beh of PGnet_1 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity carry_select_N4_7 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_N4_7;

architecture SYN_beh of carry_select_N4_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_generic_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_13
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_14
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sel, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, net2289, net2290 :
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_GEN_NBIT4_14 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => net2290);
   RCA2 : RCA_GEN_NBIT4_13 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => net2289);
   MUX1 : mux21_generic_NBIT4_7 port map( A(3) => S0_3_port, A(2) => S0_2_port,
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => sel, Y(3) => S(3), Y(2) =>
                           S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : INV_X1 port map( A => Cin, ZN => sel);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity carry_select_N4_6 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_N4_6;

architecture SYN_beh of carry_select_N4_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_generic_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_11
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_12
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sel, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, net2289, net2290 :
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_GEN_NBIT4_12 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => net2290);
   RCA2 : RCA_GEN_NBIT4_11 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => net2289);
   MUX1 : mux21_generic_NBIT4_6 port map( A(3) => S0_3_port, A(2) => S0_2_port,
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => sel, Y(3) => S(3), Y(2) =>
                           S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : INV_X1 port map( A => Cin, ZN => sel);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity carry_select_N4_5 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_N4_5;

architecture SYN_beh of carry_select_N4_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_generic_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_9
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_10
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sel, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, net2289, net2290 :
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_GEN_NBIT4_10 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => net2290);
   RCA2 : RCA_GEN_NBIT4_9 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => net2289);
   MUX1 : mux21_generic_NBIT4_5 port map( A(3) => S0_3_port, A(2) => S0_2_port,
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => sel, Y(3) => S(3), Y(2) =>
                           S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : INV_X1 port map( A => Cin, ZN => sel);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity carry_select_N4_4 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_N4_4;

architecture SYN_beh of carry_select_N4_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_generic_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_7
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_8
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sel, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, net2289, net2290 :
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_GEN_NBIT4_8 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => net2290);
   RCA2 : RCA_GEN_NBIT4_7 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => net2289);
   MUX1 : mux21_generic_NBIT4_4 port map( A(3) => S0_3_port, A(2) => S0_2_port,
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => sel, Y(3) => S(3), Y(2) =>
                           S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : INV_X1 port map( A => Cin, ZN => sel);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity carry_select_N4_3 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_N4_3;

architecture SYN_beh of carry_select_N4_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_generic_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_5
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_6
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sel, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, net2289, net2290 :
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_GEN_NBIT4_6 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => net2290);
   RCA2 : RCA_GEN_NBIT4_5 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => net2289);
   MUX1 : mux21_generic_NBIT4_3 port map( A(3) => S0_3_port, A(2) => S0_2_port,
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => sel, Y(3) => S(3), Y(2) =>
                           S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : INV_X1 port map( A => Cin, ZN => sel);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity carry_select_N4_2 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_N4_2;

architecture SYN_beh of carry_select_N4_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_generic_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_3
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_4
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sel, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, net2289, net2290 :
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_GEN_NBIT4_4 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => net2290);
   RCA2 : RCA_GEN_NBIT4_3 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => net2289);
   MUX1 : mux21_generic_NBIT4_2 port map( A(3) => S0_3_port, A(2) => S0_2_port,
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => sel, Y(3) => S(3), Y(2) =>
                           S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : INV_X1 port map( A => Cin, ZN => sel);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity carry_select_N4_1 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_N4_1;

architecture SYN_beh of carry_select_N4_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_generic_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_1
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_2
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sel, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, net2289, net2290 :
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_GEN_NBIT4_2 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => net2290);
   RCA2 : RCA_GEN_NBIT4_1 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => net2289);
   MUX1 : mux21_generic_NBIT4_1 port map( A(3) => S0_3_port, A(2) => S0_2_port,
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => sel, Y(3) => S(3), Y(2) =>
                           S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : INV_X1 port map( A => Cin, ZN => sel);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_43 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_43;

architecture SYN_beh of PG_43 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_42 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_42;

architecture SYN_beh of PG_42 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_41 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_41;

architecture SYN_beh of PG_41 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_40 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_40;

architecture SYN_beh of PG_40 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_39 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_39;

architecture SYN_beh of PG_39 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_38 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_38;

architecture SYN_beh of PG_38 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_37 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_37;

architecture SYN_beh of PG_37 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_36 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_36;

architecture SYN_beh of PG_36 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_35 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_35;

architecture SYN_beh of PG_35 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_34 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_34;

architecture SYN_beh of PG_34 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_33 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_33;

architecture SYN_beh of PG_33 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_32 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_32;

architecture SYN_beh of PG_32 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_31 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_31;

architecture SYN_beh of PG_31 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_30 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_30;

architecture SYN_beh of PG_30 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_29 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_29;

architecture SYN_beh of PG_29 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_28 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_28;

architecture SYN_beh of PG_28 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_27 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_27;

architecture SYN_beh of PG_27 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_26 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_26;

architecture SYN_beh of PG_26 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_25 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_25;

architecture SYN_beh of PG_25 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_24 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_24;

architecture SYN_beh of PG_24 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_23 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_23;

architecture SYN_beh of PG_23 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_22 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_22;

architecture SYN_beh of PG_22 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_21 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_21;

architecture SYN_beh of PG_21 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_20 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_20;

architecture SYN_beh of PG_20 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_19 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_19;

architecture SYN_beh of PG_19 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_18 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_18;

architecture SYN_beh of PG_18 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_17 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_17;

architecture SYN_beh of PG_17 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_16 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_16;

architecture SYN_beh of PG_16 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_15 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_15;

architecture SYN_beh of PG_15 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_14 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_14;

architecture SYN_beh of PG_14 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_13 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_13;

architecture SYN_beh of PG_13 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_12 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_12;

architecture SYN_beh of PG_12 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_11 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_11;

architecture SYN_beh of PG_11 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_10 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_10;

architecture SYN_beh of PG_10 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_9 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_9;

architecture SYN_beh of PG_9 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_8 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_8;

architecture SYN_beh of PG_8 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_7 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_7;

architecture SYN_beh of PG_7 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_6 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_6;

architecture SYN_beh of PG_6 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_5 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_5;

architecture SYN_beh of PG_5 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_4 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_4;

architecture SYN_beh of PG_4 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_3 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_3;

architecture SYN_beh of PG_3 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_2 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_2;

architecture SYN_beh of PG_2 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_1 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_1;

architecture SYN_beh of PG_1 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sparse_tree_carry_gen_4bits_7 is

   port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, G :
         out std_logic);

end sparse_tree_carry_gen_4bits_7;

architecture SYN_beh of sparse_tree_carry_gen_4bits_7 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component PG_19
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_20
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_21
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_19
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_20
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_21
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   signal X_Logic0_port, P0_3_port, P0_2_port, P0_1_port, P0_0_port, G0_3_port,
      G0_2_port, G0_1_port, G0_0_port, G1_1_port, G1_0_port, P1_1_port, 
      P1_0_port, n1, n2, n3 : std_logic;

begin
   
   X_Logic0_port <= '0';
   pg1_1 : PGnet_21 port map( A => A(1), B => B(1), C => X_Logic0_port, P => 
                           P0_1_port, G => G0_1_port);
   pg1_2 : PGnet_20 port map( A => A(2), B => B(2), C => X_Logic0_port, P => 
                           P0_2_port, G => G0_2_port);
   pg1_3 : PGnet_19 port map( A => A(3), B => B(3), C => X_Logic0_port, P => 
                           P0_3_port, G => G0_3_port);
   pg2_0 : PG_21 port map( A => P0_1_port, B => P0_0_port, C => G0_1_port, D =>
                           G0_0_port, P => P1_0_port, G => G1_0_port);
   pg2_1 : PG_20 port map( A => P0_3_port, B => P0_2_port, C => G0_3_port, D =>
                           G0_2_port, P => P1_1_port, G => G1_1_port);
   pgg : PG_19 port map( A => P1_1_port, B => P1_0_port, C => G1_1_port, D => 
                           G1_0_port, P => P, G => G);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => P0_0_port);
   U3 : INV_X1 port map( A => n1, ZN => G0_0_port);
   U4 : AOI21_X1 port map( B1 => B(0), B2 => A(0), A => n2, ZN => n1);
   U5 : INV_X1 port map( A => n3, ZN => n2);
   U6 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => c_in, ZN => n3);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sparse_tree_carry_gen_4bits_6 is

   port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, G :
         out std_logic);

end sparse_tree_carry_gen_4bits_6;

architecture SYN_beh of sparse_tree_carry_gen_4bits_6 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component PG_16
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_17
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_18
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_16
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_17
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_18
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   signal X_Logic0_port, P0_3_port, P0_2_port, P0_1_port, P0_0_port, G0_3_port,
      G0_2_port, G0_1_port, G0_0_port, G1_1_port, G1_0_port, P1_1_port, 
      P1_0_port, n1, n2, n3 : std_logic;

begin
   
   X_Logic0_port <= '0';
   pg1_1 : PGnet_18 port map( A => A(1), B => B(1), C => X_Logic0_port, P => 
                           P0_1_port, G => G0_1_port);
   pg1_2 : PGnet_17 port map( A => A(2), B => B(2), C => X_Logic0_port, P => 
                           P0_2_port, G => G0_2_port);
   pg1_3 : PGnet_16 port map( A => A(3), B => B(3), C => X_Logic0_port, P => 
                           P0_3_port, G => G0_3_port);
   pg2_0 : PG_18 port map( A => P0_1_port, B => P0_0_port, C => G0_1_port, D =>
                           G0_0_port, P => P1_0_port, G => G1_0_port);
   pg2_1 : PG_17 port map( A => P0_3_port, B => P0_2_port, C => G0_3_port, D =>
                           G0_2_port, P => P1_1_port, G => G1_1_port);
   pgg : PG_16 port map( A => P1_1_port, B => P1_0_port, C => G1_1_port, D => 
                           G1_0_port, P => P, G => G);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => P0_0_port);
   U3 : INV_X1 port map( A => n1, ZN => G0_0_port);
   U4 : AOI21_X1 port map( B1 => B(0), B2 => A(0), A => n2, ZN => n1);
   U5 : INV_X1 port map( A => n3, ZN => n2);
   U6 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => c_in, ZN => n3);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sparse_tree_carry_gen_4bits_5 is

   port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, G :
         out std_logic);

end sparse_tree_carry_gen_4bits_5;

architecture SYN_beh of sparse_tree_carry_gen_4bits_5 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component PG_13
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_14
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_15
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_13
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_14
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_15
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   signal X_Logic0_port, P0_3_port, P0_2_port, P0_1_port, P0_0_port, G0_3_port,
      G0_2_port, G0_1_port, G0_0_port, G1_1_port, G1_0_port, P1_1_port, 
      P1_0_port, n1, n2, n3 : std_logic;

begin
   
   X_Logic0_port <= '0';
   pg1_1 : PGnet_15 port map( A => A(1), B => B(1), C => X_Logic0_port, P => 
                           P0_1_port, G => G0_1_port);
   pg1_2 : PGnet_14 port map( A => A(2), B => B(2), C => X_Logic0_port, P => 
                           P0_2_port, G => G0_2_port);
   pg1_3 : PGnet_13 port map( A => A(3), B => B(3), C => X_Logic0_port, P => 
                           P0_3_port, G => G0_3_port);
   pg2_0 : PG_15 port map( A => P0_1_port, B => P0_0_port, C => G0_1_port, D =>
                           G0_0_port, P => P1_0_port, G => G1_0_port);
   pg2_1 : PG_14 port map( A => P0_3_port, B => P0_2_port, C => G0_3_port, D =>
                           G0_2_port, P => P1_1_port, G => G1_1_port);
   pgg : PG_13 port map( A => P1_1_port, B => P1_0_port, C => G1_1_port, D => 
                           G1_0_port, P => P, G => G);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => P0_0_port);
   U3 : INV_X1 port map( A => n1, ZN => G0_0_port);
   U4 : AOI21_X1 port map( B1 => B(0), B2 => A(0), A => n2, ZN => n1);
   U5 : INV_X1 port map( A => n3, ZN => n2);
   U6 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => c_in, ZN => n3);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sparse_tree_carry_gen_4bits_4 is

   port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, G :
         out std_logic);

end sparse_tree_carry_gen_4bits_4;

architecture SYN_beh of sparse_tree_carry_gen_4bits_4 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component PG_10
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_11
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_12
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_10
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_11
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_12
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   signal X_Logic0_port, P0_3_port, P0_2_port, P0_1_port, P0_0_port, G0_3_port,
      G0_2_port, G0_1_port, G0_0_port, G1_1_port, G1_0_port, P1_1_port, 
      P1_0_port, n1, n2, n3 : std_logic;

begin
   
   X_Logic0_port <= '0';
   pg1_1 : PGnet_12 port map( A => A(1), B => B(1), C => X_Logic0_port, P => 
                           P0_1_port, G => G0_1_port);
   pg1_2 : PGnet_11 port map( A => A(2), B => B(2), C => X_Logic0_port, P => 
                           P0_2_port, G => G0_2_port);
   pg1_3 : PGnet_10 port map( A => A(3), B => B(3), C => X_Logic0_port, P => 
                           P0_3_port, G => G0_3_port);
   pg2_0 : PG_12 port map( A => P0_1_port, B => P0_0_port, C => G0_1_port, D =>
                           G0_0_port, P => P1_0_port, G => G1_0_port);
   pg2_1 : PG_11 port map( A => P0_3_port, B => P0_2_port, C => G0_3_port, D =>
                           G0_2_port, P => P1_1_port, G => G1_1_port);
   pgg : PG_10 port map( A => P1_1_port, B => P1_0_port, C => G1_1_port, D => 
                           G1_0_port, P => P, G => G);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => P0_0_port);
   U3 : INV_X1 port map( A => n1, ZN => G0_0_port);
   U4 : AOI21_X1 port map( B1 => B(0), B2 => A(0), A => n2, ZN => n1);
   U5 : INV_X1 port map( A => n3, ZN => n2);
   U6 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => c_in, ZN => n3);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sparse_tree_carry_gen_4bits_3 is

   port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, G :
         out std_logic);

end sparse_tree_carry_gen_4bits_3;

architecture SYN_beh of sparse_tree_carry_gen_4bits_3 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component PG_7
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_8
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_9
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_7
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_8
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_9
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   signal X_Logic0_port, P0_3_port, P0_2_port, P0_1_port, P0_0_port, G0_3_port,
      G0_2_port, G0_1_port, G0_0_port, G1_1_port, G1_0_port, P1_1_port, 
      P1_0_port, n1, n2, n3 : std_logic;

begin
   
   X_Logic0_port <= '0';
   pg1_1 : PGnet_9 port map( A => A(1), B => B(1), C => X_Logic0_port, P => 
                           P0_1_port, G => G0_1_port);
   pg1_2 : PGnet_8 port map( A => A(2), B => B(2), C => X_Logic0_port, P => 
                           P0_2_port, G => G0_2_port);
   pg1_3 : PGnet_7 port map( A => A(3), B => B(3), C => X_Logic0_port, P => 
                           P0_3_port, G => G0_3_port);
   pg2_0 : PG_9 port map( A => P0_1_port, B => P0_0_port, C => G0_1_port, D => 
                           G0_0_port, P => P1_0_port, G => G1_0_port);
   pg2_1 : PG_8 port map( A => P0_3_port, B => P0_2_port, C => G0_3_port, D => 
                           G0_2_port, P => P1_1_port, G => G1_1_port);
   pgg : PG_7 port map( A => P1_1_port, B => P1_0_port, C => G1_1_port, D => 
                           G1_0_port, P => P, G => G);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => P0_0_port);
   U3 : INV_X1 port map( A => n1, ZN => G0_0_port);
   U4 : AOI21_X1 port map( B1 => B(0), B2 => A(0), A => n2, ZN => n1);
   U5 : INV_X1 port map( A => n3, ZN => n2);
   U6 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => c_in, ZN => n3);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sparse_tree_carry_gen_4bits_2 is

   port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, G :
         out std_logic);

end sparse_tree_carry_gen_4bits_2;

architecture SYN_beh of sparse_tree_carry_gen_4bits_2 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component PG_4
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_5
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_6
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_4
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_5
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_6
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   signal X_Logic0_port, P0_3_port, P0_2_port, P0_1_port, P0_0_port, G0_3_port,
      G0_2_port, G0_1_port, G0_0_port, G1_1_port, G1_0_port, P1_1_port, 
      P1_0_port, n1, n2, n3 : std_logic;

begin
   
   X_Logic0_port <= '0';
   pg1_1 : PGnet_6 port map( A => A(1), B => B(1), C => X_Logic0_port, P => 
                           P0_1_port, G => G0_1_port);
   pg1_2 : PGnet_5 port map( A => A(2), B => B(2), C => X_Logic0_port, P => 
                           P0_2_port, G => G0_2_port);
   pg1_3 : PGnet_4 port map( A => A(3), B => B(3), C => X_Logic0_port, P => 
                           P0_3_port, G => G0_3_port);
   pg2_0 : PG_6 port map( A => P0_1_port, B => P0_0_port, C => G0_1_port, D => 
                           G0_0_port, P => P1_0_port, G => G1_0_port);
   pg2_1 : PG_5 port map( A => P0_3_port, B => P0_2_port, C => G0_3_port, D => 
                           G0_2_port, P => P1_1_port, G => G1_1_port);
   pgg : PG_4 port map( A => P1_1_port, B => P1_0_port, C => G1_1_port, D => 
                           G1_0_port, P => P, G => G);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => P0_0_port);
   U3 : INV_X1 port map( A => n1, ZN => G0_0_port);
   U4 : AOI21_X1 port map( B1 => B(0), B2 => A(0), A => n2, ZN => n1);
   U5 : INV_X1 port map( A => n3, ZN => n2);
   U6 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => c_in, ZN => n3);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sparse_tree_carry_gen_4bits_1 is

   port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, G :
         out std_logic);

end sparse_tree_carry_gen_4bits_1;

architecture SYN_beh of sparse_tree_carry_gen_4bits_1 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component PG_1
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_2
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_3
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_1
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_2
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_3
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   signal X_Logic0_port, P0_3_port, P0_2_port, P0_1_port, P0_0_port, G0_3_port,
      G0_2_port, G0_1_port, G0_0_port, G1_1_port, G1_0_port, P1_1_port, 
      P1_0_port, n1, n2, n3 : std_logic;

begin
   
   X_Logic0_port <= '0';
   pg1_1 : PGnet_3 port map( A => A(1), B => B(1), C => X_Logic0_port, P => 
                           P0_1_port, G => G0_1_port);
   pg1_2 : PGnet_2 port map( A => A(2), B => B(2), C => X_Logic0_port, P => 
                           P0_2_port, G => G0_2_port);
   pg1_3 : PGnet_1 port map( A => A(3), B => B(3), C => X_Logic0_port, P => 
                           P0_3_port, G => G0_3_port);
   pg2_0 : PG_3 port map( A => P0_1_port, B => P0_0_port, C => G0_1_port, D => 
                           G0_0_port, P => P1_0_port, G => G1_0_port);
   pg2_1 : PG_2 port map( A => P0_3_port, B => P0_2_port, C => G0_3_port, D => 
                           G0_2_port, P => P1_1_port, G => G1_1_port);
   pgg : PG_1 port map( A => P1_1_port, B => P1_0_port, C => G1_1_port, D => 
                           G1_0_port, P => P, G => G);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => P0_0_port);
   U3 : INV_X1 port map( A => n1, ZN => G0_0_port);
   U4 : AOI21_X1 port map( B1 => B(0), B2 => A(0), A => n2, ZN => n1);
   U5 : INV_X1 port map( A => n3, ZN => n2);
   U6 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => c_in, ZN => n3);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_95 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_95;

architecture SYN_BEHAVIORAL of FA_95 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_94 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_94;

architecture SYN_BEHAVIORAL of FA_94 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_93 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_93;

architecture SYN_BEHAVIORAL of FA_93 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_92 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_92;

architecture SYN_BEHAVIORAL of FA_92 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_91 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_91;

architecture SYN_BEHAVIORAL of FA_91 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_90 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_90;

architecture SYN_BEHAVIORAL of FA_90 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_89 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_89;

architecture SYN_BEHAVIORAL of FA_89 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_88 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_88;

architecture SYN_BEHAVIORAL of FA_88 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_87 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_87;

architecture SYN_BEHAVIORAL of FA_87 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_86 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_86;

architecture SYN_BEHAVIORAL of FA_86 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_85 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_85;

architecture SYN_BEHAVIORAL of FA_85 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_84 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_84;

architecture SYN_BEHAVIORAL of FA_84 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_83 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_83;

architecture SYN_BEHAVIORAL of FA_83 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_82 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_82;

architecture SYN_BEHAVIORAL of FA_82 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_81 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_81;

architecture SYN_BEHAVIORAL of FA_81 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_80 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_80;

architecture SYN_BEHAVIORAL of FA_80 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_79 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_79;

architecture SYN_BEHAVIORAL of FA_79 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_78 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_78;

architecture SYN_BEHAVIORAL of FA_78 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_77 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_77;

architecture SYN_BEHAVIORAL of FA_77 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_76 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_76;

architecture SYN_BEHAVIORAL of FA_76 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_75 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_75;

architecture SYN_BEHAVIORAL of FA_75 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_74 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_74;

architecture SYN_BEHAVIORAL of FA_74 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_73 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_73;

architecture SYN_BEHAVIORAL of FA_73 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_72 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_72;

architecture SYN_BEHAVIORAL of FA_72 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_71 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_71;

architecture SYN_BEHAVIORAL of FA_71 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_70 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_70;

architecture SYN_BEHAVIORAL of FA_70 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_69 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_69;

architecture SYN_BEHAVIORAL of FA_69 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_68 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_68;

architecture SYN_BEHAVIORAL of FA_68 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_67 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_67;

architecture SYN_BEHAVIORAL of FA_67 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_66 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_66;

architecture SYN_BEHAVIORAL of FA_66 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_65 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_65;

architecture SYN_BEHAVIORAL of FA_65 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_64 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_64;

architecture SYN_BEHAVIORAL of FA_64 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL_architecture of FA_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL_architecture2 of FA_58 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL_architecture3 of FA_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL_architecture of FA_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL_architecture2 of FA_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL_architecture3 of FA_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL_architecture of FA_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL_architecture2 of FA_50 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL_architecture3 of FA_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL_architecture of FA_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL_architecture2 of FA_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL_architecture3 of FA_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL_architecture of FA_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL_architecture2 of FA_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL_architecture3 of FA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL_architecture of FA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL_architecture2 of FA_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL_architecture3 of FA_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL_architecture of FA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL_architecture2 of FA_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL_architecture3 of FA_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL_architecture of FA_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL_architecture2 of FA_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL_architecture3 of FA_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL_architecture of FA_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL_architecture2 of FA_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL_architecture3 of FA_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL_architecture of FA_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL_architecture2 of FA_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL_architecture3 of FA_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL_architecture of FA_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL_architecture2 of FA_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL_architecture3 of FA_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL_architecture of FA_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL_architecture2 of FA_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL_architecture3 of FA_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL_architecture of FA_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL_architecture2 of FA_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL_architecture3 of FA_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL_architecture of FA_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL_architecture2 of FA_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL_architecture3 of FA_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL_architecture of FA_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL_architecture2 of FA_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture2;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL_architecture3 of FA_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL_architecture3;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N5_2 is

   port( data : in std_logic_vector (4 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (4 downto 0));

end registro_N5_2;

architecture SYN_behaviour of registro_N5_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n1, n2, n3, n4, n5,
      net43512, net43513, net43514, net43515, net43516 : std_logic;

begin
   Q <= ( Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_4_inst : DFFR_X1 port map( D => n1, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43516);
   Q_reg_3_inst : DFFR_X1 port map( D => n2, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43515);
   Q_reg_2_inst : DFFR_X1 port map( D => n3, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43514);
   Q_reg_1_inst : DFFR_X1 port map( D => n4, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43513);
   Q_reg_0_inst : DFFR_X1 port map( D => n5, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43512);
   U2 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n1);
   U3 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n2);
   U4 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n3);
   U5 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n4);
   U6 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n5);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N5_1 is

   port( data : in std_logic_vector (4 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (4 downto 0));

end registro_N5_1;

architecture SYN_behaviour of registro_N5_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n1, n2, n3, n4, n5,
      net43507, net43508, net43509, net43510, net43511 : std_logic;

begin
   Q <= ( Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_4_inst : DFFR_X1 port map( D => n1, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43511);
   Q_reg_3_inst : DFFR_X1 port map( D => n2, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43510);
   Q_reg_2_inst : DFFR_X1 port map( D => n3, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43509);
   Q_reg_1_inst : DFFR_X1 port map( D => n4, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43508);
   Q_reg_0_inst : DFFR_X1 port map( D => n5, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43507);
   U2 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n1);
   U3 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n2);
   U4 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n3);
   U5 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n4);
   U6 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n5);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N32_8 is

   port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end registro_N32_8;

architecture SYN_behaviour of registro_N32_8 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , net43475, net43476, net43477, net43478, net43479, net43480, net43481, 
      net43482, net43483, net43484, net43485, net43486, net43487, net43488, 
      net43489, net43490, net43491, net43492, net43493, net43494, net43495, 
      net43496, net43497, net43498, net43499, net43500, net43501, net43502, 
      net43503, net43504, net43505, net43506 : std_logic;

begin
   Q <= ( Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => clock, RN => clear, Q => 
                           Q_31_port, QN => net43506);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => clock, RN => clear, Q => 
                           Q_30_port, QN => net43505);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => clock, RN => clear, Q => 
                           Q_29_port, QN => net43504);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => clock, RN => clear, Q => 
                           Q_28_port, QN => net43503);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => clock, RN => clear, Q => 
                           Q_27_port, QN => net43502);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => clock, RN => clear, Q => 
                           Q_26_port, QN => net43501);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => clock, RN => clear, Q => 
                           Q_25_port, QN => net43500);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => clock, RN => clear, Q => 
                           Q_24_port, QN => net43499);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => clock, RN => clear, Q => 
                           Q_23_port, QN => net43498);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => clock, RN => clear, Q => 
                           Q_22_port, QN => net43497);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => clock, RN => clear, Q => 
                           Q_21_port, QN => net43496);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => clock, RN => clear, Q => 
                           Q_20_port, QN => net43495);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => clock, RN => clear, Q => 
                           Q_19_port, QN => net43494);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => clock, RN => clear, Q => 
                           Q_18_port, QN => net43493);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => clock, RN => clear, Q => 
                           Q_17_port, QN => net43492);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => clock, RN => clear, Q => 
                           Q_16_port, QN => net43491);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => clock, RN => clear, Q => 
                           Q_15_port, QN => net43490);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => clock, RN => clear, Q => 
                           Q_14_port, QN => net43489);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => clock, RN => clear, Q => 
                           Q_13_port, QN => net43488);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => clock, RN => clear, Q => 
                           Q_12_port, QN => net43487);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => clock, RN => clear, Q => 
                           Q_11_port, QN => net43486);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => clock, RN => clear, Q => 
                           Q_10_port, QN => net43485);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => clock, RN => clear, Q => 
                           Q_9_port, QN => net43484);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => clock, RN => clear, Q => 
                           Q_8_port, QN => net43483);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => clock, RN => clear, Q => 
                           Q_7_port, QN => net43482);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => clock, RN => clear, Q => 
                           Q_6_port, QN => net43481);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => clock, RN => clear, Q => 
                           Q_5_port, QN => net43480);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43479);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43478);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43477);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43476);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43475);
   U2 : MUX2_X1 port map( A => Q_31_port, B => data(31), S => enable, Z => n1);
   U3 : MUX2_X1 port map( A => Q_30_port, B => data(30), S => enable, Z => n2);
   U4 : MUX2_X1 port map( A => Q_29_port, B => data(29), S => enable, Z => n3);
   U5 : MUX2_X1 port map( A => Q_28_port, B => data(28), S => enable, Z => n4);
   U6 : MUX2_X1 port map( A => Q_27_port, B => data(27), S => enable, Z => n5);
   U7 : MUX2_X1 port map( A => Q_26_port, B => data(26), S => enable, Z => n6);
   U8 : MUX2_X1 port map( A => Q_25_port, B => data(25), S => enable, Z => n7);
   U9 : MUX2_X1 port map( A => Q_24_port, B => data(24), S => enable, Z => n8);
   U10 : MUX2_X1 port map( A => Q_23_port, B => data(23), S => enable, Z => n9)
                           ;
   U11 : MUX2_X1 port map( A => Q_22_port, B => data(22), S => enable, Z => n10
                           );
   U12 : MUX2_X1 port map( A => Q_21_port, B => data(21), S => enable, Z => n11
                           );
   U13 : MUX2_X1 port map( A => Q_20_port, B => data(20), S => enable, Z => n12
                           );
   U14 : MUX2_X1 port map( A => Q_19_port, B => data(19), S => enable, Z => n13
                           );
   U15 : MUX2_X1 port map( A => Q_18_port, B => data(18), S => enable, Z => n14
                           );
   U16 : MUX2_X1 port map( A => Q_17_port, B => data(17), S => enable, Z => n15
                           );
   U17 : MUX2_X1 port map( A => Q_16_port, B => data(16), S => enable, Z => n16
                           );
   U18 : MUX2_X1 port map( A => Q_15_port, B => data(15), S => enable, Z => n17
                           );
   U19 : MUX2_X1 port map( A => Q_14_port, B => data(14), S => enable, Z => n18
                           );
   U20 : MUX2_X1 port map( A => Q_13_port, B => data(13), S => enable, Z => n19
                           );
   U21 : MUX2_X1 port map( A => Q_12_port, B => data(12), S => enable, Z => n20
                           );
   U22 : MUX2_X1 port map( A => Q_11_port, B => data(11), S => enable, Z => n21
                           );
   U23 : MUX2_X1 port map( A => Q_10_port, B => data(10), S => enable, Z => n22
                           );
   U24 : MUX2_X1 port map( A => Q_9_port, B => data(9), S => enable, Z => n23);
   U25 : MUX2_X1 port map( A => Q_8_port, B => data(8), S => enable, Z => n24);
   U26 : MUX2_X1 port map( A => Q_7_port, B => data(7), S => enable, Z => n25);
   U27 : MUX2_X1 port map( A => Q_6_port, B => data(6), S => enable, Z => n26);
   U28 : MUX2_X1 port map( A => Q_5_port, B => data(5), S => enable, Z => n27);
   U29 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n28);
   U30 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n29);
   U31 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n30);
   U32 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n31);
   U33 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n32);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N32_7 is

   port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end registro_N32_7;

architecture SYN_behaviour of registro_N32_7 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , net43443, net43444, net43445, net43446, net43447, net43448, net43449, 
      net43450, net43451, net43452, net43453, net43454, net43455, net43456, 
      net43457, net43458, net43459, net43460, net43461, net43462, net43463, 
      net43464, net43465, net43466, net43467, net43468, net43469, net43470, 
      net43471, net43472, net43473, net43474 : std_logic;

begin
   Q <= ( Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => clock, RN => clear, Q => 
                           Q_31_port, QN => net43474);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => clock, RN => clear, Q => 
                           Q_30_port, QN => net43473);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => clock, RN => clear, Q => 
                           Q_29_port, QN => net43472);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => clock, RN => clear, Q => 
                           Q_28_port, QN => net43471);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => clock, RN => clear, Q => 
                           Q_27_port, QN => net43470);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => clock, RN => clear, Q => 
                           Q_26_port, QN => net43469);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => clock, RN => clear, Q => 
                           Q_25_port, QN => net43468);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => clock, RN => clear, Q => 
                           Q_24_port, QN => net43467);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => clock, RN => clear, Q => 
                           Q_23_port, QN => net43466);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => clock, RN => clear, Q => 
                           Q_22_port, QN => net43465);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => clock, RN => clear, Q => 
                           Q_21_port, QN => net43464);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => clock, RN => clear, Q => 
                           Q_20_port, QN => net43463);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => clock, RN => clear, Q => 
                           Q_19_port, QN => net43462);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => clock, RN => clear, Q => 
                           Q_18_port, QN => net43461);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => clock, RN => clear, Q => 
                           Q_17_port, QN => net43460);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => clock, RN => clear, Q => 
                           Q_16_port, QN => net43459);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => clock, RN => clear, Q => 
                           Q_15_port, QN => net43458);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => clock, RN => clear, Q => 
                           Q_14_port, QN => net43457);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => clock, RN => clear, Q => 
                           Q_13_port, QN => net43456);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => clock, RN => clear, Q => 
                           Q_12_port, QN => net43455);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => clock, RN => clear, Q => 
                           Q_11_port, QN => net43454);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => clock, RN => clear, Q => 
                           Q_10_port, QN => net43453);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => clock, RN => clear, Q => 
                           Q_9_port, QN => net43452);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => clock, RN => clear, Q => 
                           Q_8_port, QN => net43451);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => clock, RN => clear, Q => 
                           Q_7_port, QN => net43450);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => clock, RN => clear, Q => 
                           Q_6_port, QN => net43449);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => clock, RN => clear, Q => 
                           Q_5_port, QN => net43448);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43447);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43446);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43445);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43444);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43443);
   U2 : MUX2_X1 port map( A => Q_31_port, B => data(31), S => enable, Z => n1);
   U3 : MUX2_X1 port map( A => Q_30_port, B => data(30), S => enable, Z => n2);
   U4 : MUX2_X1 port map( A => Q_29_port, B => data(29), S => enable, Z => n3);
   U5 : MUX2_X1 port map( A => Q_28_port, B => data(28), S => enable, Z => n4);
   U6 : MUX2_X1 port map( A => Q_27_port, B => data(27), S => enable, Z => n5);
   U7 : MUX2_X1 port map( A => Q_26_port, B => data(26), S => enable, Z => n6);
   U8 : MUX2_X1 port map( A => Q_25_port, B => data(25), S => enable, Z => n7);
   U9 : MUX2_X1 port map( A => Q_24_port, B => data(24), S => enable, Z => n8);
   U10 : MUX2_X1 port map( A => Q_23_port, B => data(23), S => enable, Z => n9)
                           ;
   U11 : MUX2_X1 port map( A => Q_22_port, B => data(22), S => enable, Z => n10
                           );
   U12 : MUX2_X1 port map( A => Q_21_port, B => data(21), S => enable, Z => n11
                           );
   U13 : MUX2_X1 port map( A => Q_20_port, B => data(20), S => enable, Z => n12
                           );
   U14 : MUX2_X1 port map( A => Q_19_port, B => data(19), S => enable, Z => n13
                           );
   U15 : MUX2_X1 port map( A => Q_18_port, B => data(18), S => enable, Z => n14
                           );
   U16 : MUX2_X1 port map( A => Q_17_port, B => data(17), S => enable, Z => n15
                           );
   U17 : MUX2_X1 port map( A => Q_16_port, B => data(16), S => enable, Z => n16
                           );
   U18 : MUX2_X1 port map( A => Q_15_port, B => data(15), S => enable, Z => n17
                           );
   U19 : MUX2_X1 port map( A => Q_14_port, B => data(14), S => enable, Z => n18
                           );
   U20 : MUX2_X1 port map( A => Q_13_port, B => data(13), S => enable, Z => n19
                           );
   U21 : MUX2_X1 port map( A => Q_12_port, B => data(12), S => enable, Z => n20
                           );
   U22 : MUX2_X1 port map( A => Q_11_port, B => data(11), S => enable, Z => n21
                           );
   U23 : MUX2_X1 port map( A => Q_10_port, B => data(10), S => enable, Z => n22
                           );
   U24 : MUX2_X1 port map( A => Q_9_port, B => data(9), S => enable, Z => n23);
   U25 : MUX2_X1 port map( A => Q_8_port, B => data(8), S => enable, Z => n24);
   U26 : MUX2_X1 port map( A => Q_7_port, B => data(7), S => enable, Z => n25);
   U27 : MUX2_X1 port map( A => Q_6_port, B => data(6), S => enable, Z => n26);
   U28 : MUX2_X1 port map( A => Q_5_port, B => data(5), S => enable, Z => n27);
   U29 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n28);
   U30 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n29);
   U31 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n30);
   U32 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n31);
   U33 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n32);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N32_6 is

   port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end registro_N32_6;

architecture SYN_behaviour of registro_N32_6 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , net43411, net43412, net43413, net43414, net43415, net43416, net43417, 
      net43418, net43419, net43420, net43421, net43422, net43423, net43424, 
      net43425, net43426, net43427, net43428, net43429, net43430, net43431, 
      net43432, net43433, net43434, net43435, net43436, net43437, net43438, 
      net43439, net43440, net43441, net43442 : std_logic;

begin
   Q <= ( Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => clock, RN => clear, Q => 
                           Q_31_port, QN => net43442);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => clock, RN => clear, Q => 
                           Q_30_port, QN => net43441);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => clock, RN => clear, Q => 
                           Q_29_port, QN => net43440);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => clock, RN => clear, Q => 
                           Q_28_port, QN => net43439);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => clock, RN => clear, Q => 
                           Q_27_port, QN => net43438);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => clock, RN => clear, Q => 
                           Q_26_port, QN => net43437);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => clock, RN => clear, Q => 
                           Q_25_port, QN => net43436);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => clock, RN => clear, Q => 
                           Q_24_port, QN => net43435);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => clock, RN => clear, Q => 
                           Q_23_port, QN => net43434);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => clock, RN => clear, Q => 
                           Q_22_port, QN => net43433);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => clock, RN => clear, Q => 
                           Q_21_port, QN => net43432);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => clock, RN => clear, Q => 
                           Q_20_port, QN => net43431);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => clock, RN => clear, Q => 
                           Q_19_port, QN => net43430);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => clock, RN => clear, Q => 
                           Q_18_port, QN => net43429);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => clock, RN => clear, Q => 
                           Q_17_port, QN => net43428);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => clock, RN => clear, Q => 
                           Q_16_port, QN => net43427);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => clock, RN => clear, Q => 
                           Q_15_port, QN => net43426);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => clock, RN => clear, Q => 
                           Q_14_port, QN => net43425);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => clock, RN => clear, Q => 
                           Q_13_port, QN => net43424);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => clock, RN => clear, Q => 
                           Q_12_port, QN => net43423);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => clock, RN => clear, Q => 
                           Q_11_port, QN => net43422);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => clock, RN => clear, Q => 
                           Q_10_port, QN => net43421);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => clock, RN => clear, Q => 
                           Q_9_port, QN => net43420);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => clock, RN => clear, Q => 
                           Q_8_port, QN => net43419);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => clock, RN => clear, Q => 
                           Q_7_port, QN => net43418);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => clock, RN => clear, Q => 
                           Q_6_port, QN => net43417);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => clock, RN => clear, Q => 
                           Q_5_port, QN => net43416);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43415);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43414);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43413);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43412);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43411);
   U2 : MUX2_X1 port map( A => Q_31_port, B => data(31), S => enable, Z => n1);
   U3 : MUX2_X1 port map( A => Q_30_port, B => data(30), S => enable, Z => n2);
   U4 : MUX2_X1 port map( A => Q_29_port, B => data(29), S => enable, Z => n3);
   U5 : MUX2_X1 port map( A => Q_28_port, B => data(28), S => enable, Z => n4);
   U6 : MUX2_X1 port map( A => Q_27_port, B => data(27), S => enable, Z => n5);
   U7 : MUX2_X1 port map( A => Q_26_port, B => data(26), S => enable, Z => n6);
   U8 : MUX2_X1 port map( A => Q_25_port, B => data(25), S => enable, Z => n7);
   U9 : MUX2_X1 port map( A => Q_24_port, B => data(24), S => enable, Z => n8);
   U10 : MUX2_X1 port map( A => Q_23_port, B => data(23), S => enable, Z => n9)
                           ;
   U11 : MUX2_X1 port map( A => Q_22_port, B => data(22), S => enable, Z => n10
                           );
   U12 : MUX2_X1 port map( A => Q_21_port, B => data(21), S => enable, Z => n11
                           );
   U13 : MUX2_X1 port map( A => Q_20_port, B => data(20), S => enable, Z => n12
                           );
   U14 : MUX2_X1 port map( A => Q_19_port, B => data(19), S => enable, Z => n13
                           );
   U15 : MUX2_X1 port map( A => Q_18_port, B => data(18), S => enable, Z => n14
                           );
   U16 : MUX2_X1 port map( A => Q_17_port, B => data(17), S => enable, Z => n15
                           );
   U17 : MUX2_X1 port map( A => Q_16_port, B => data(16), S => enable, Z => n16
                           );
   U18 : MUX2_X1 port map( A => Q_15_port, B => data(15), S => enable, Z => n17
                           );
   U19 : MUX2_X1 port map( A => Q_14_port, B => data(14), S => enable, Z => n18
                           );
   U20 : MUX2_X1 port map( A => Q_13_port, B => data(13), S => enable, Z => n19
                           );
   U21 : MUX2_X1 port map( A => Q_12_port, B => data(12), S => enable, Z => n20
                           );
   U22 : MUX2_X1 port map( A => Q_11_port, B => data(11), S => enable, Z => n21
                           );
   U23 : MUX2_X1 port map( A => Q_10_port, B => data(10), S => enable, Z => n22
                           );
   U24 : MUX2_X1 port map( A => Q_9_port, B => data(9), S => enable, Z => n23);
   U25 : MUX2_X1 port map( A => Q_8_port, B => data(8), S => enable, Z => n24);
   U26 : MUX2_X1 port map( A => Q_7_port, B => data(7), S => enable, Z => n25);
   U27 : MUX2_X1 port map( A => Q_6_port, B => data(6), S => enable, Z => n26);
   U28 : MUX2_X1 port map( A => Q_5_port, B => data(5), S => enable, Z => n27);
   U29 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n28);
   U30 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n29);
   U31 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n30);
   U32 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n31);
   U33 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n32);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N32_5 is

   port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end registro_N32_5;

architecture SYN_behaviour of registro_N32_5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , net43379, net43380, net43381, net43382, net43383, net43384, net43385, 
      net43386, net43387, net43388, net43389, net43390, net43391, net43392, 
      net43393, net43394, net43395, net43396, net43397, net43398, net43399, 
      net43400, net43401, net43402, net43403, net43404, net43405, net43406, 
      net43407, net43408, net43409, net43410 : std_logic;

begin
   Q <= ( Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => clock, RN => clear, Q => 
                           Q_31_port, QN => net43410);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => clock, RN => clear, Q => 
                           Q_30_port, QN => net43409);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => clock, RN => clear, Q => 
                           Q_29_port, QN => net43408);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => clock, RN => clear, Q => 
                           Q_28_port, QN => net43407);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => clock, RN => clear, Q => 
                           Q_27_port, QN => net43406);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => clock, RN => clear, Q => 
                           Q_26_port, QN => net43405);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => clock, RN => clear, Q => 
                           Q_25_port, QN => net43404);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => clock, RN => clear, Q => 
                           Q_24_port, QN => net43403);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => clock, RN => clear, Q => 
                           Q_23_port, QN => net43402);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => clock, RN => clear, Q => 
                           Q_22_port, QN => net43401);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => clock, RN => clear, Q => 
                           Q_21_port, QN => net43400);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => clock, RN => clear, Q => 
                           Q_20_port, QN => net43399);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => clock, RN => clear, Q => 
                           Q_19_port, QN => net43398);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => clock, RN => clear, Q => 
                           Q_18_port, QN => net43397);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => clock, RN => clear, Q => 
                           Q_17_port, QN => net43396);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => clock, RN => clear, Q => 
                           Q_16_port, QN => net43395);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => clock, RN => clear, Q => 
                           Q_15_port, QN => net43394);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => clock, RN => clear, Q => 
                           Q_14_port, QN => net43393);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => clock, RN => clear, Q => 
                           Q_13_port, QN => net43392);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => clock, RN => clear, Q => 
                           Q_12_port, QN => net43391);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => clock, RN => clear, Q => 
                           Q_11_port, QN => net43390);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => clock, RN => clear, Q => 
                           Q_10_port, QN => net43389);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => clock, RN => clear, Q => 
                           Q_9_port, QN => net43388);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => clock, RN => clear, Q => 
                           Q_8_port, QN => net43387);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => clock, RN => clear, Q => 
                           Q_7_port, QN => net43386);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => clock, RN => clear, Q => 
                           Q_6_port, QN => net43385);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => clock, RN => clear, Q => 
                           Q_5_port, QN => net43384);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43383);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43382);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43381);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43380);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43379);
   U2 : MUX2_X1 port map( A => Q_31_port, B => data(31), S => enable, Z => n1);
   U3 : MUX2_X1 port map( A => Q_30_port, B => data(30), S => enable, Z => n2);
   U4 : MUX2_X1 port map( A => Q_29_port, B => data(29), S => enable, Z => n3);
   U5 : MUX2_X1 port map( A => Q_28_port, B => data(28), S => enable, Z => n4);
   U6 : MUX2_X1 port map( A => Q_27_port, B => data(27), S => enable, Z => n5);
   U7 : MUX2_X1 port map( A => Q_26_port, B => data(26), S => enable, Z => n6);
   U8 : MUX2_X1 port map( A => Q_25_port, B => data(25), S => enable, Z => n7);
   U9 : MUX2_X1 port map( A => Q_24_port, B => data(24), S => enable, Z => n8);
   U10 : MUX2_X1 port map( A => Q_23_port, B => data(23), S => enable, Z => n9)
                           ;
   U11 : MUX2_X1 port map( A => Q_22_port, B => data(22), S => enable, Z => n10
                           );
   U12 : MUX2_X1 port map( A => Q_21_port, B => data(21), S => enable, Z => n11
                           );
   U13 : MUX2_X1 port map( A => Q_20_port, B => data(20), S => enable, Z => n12
                           );
   U14 : MUX2_X1 port map( A => Q_19_port, B => data(19), S => enable, Z => n13
                           );
   U15 : MUX2_X1 port map( A => Q_18_port, B => data(18), S => enable, Z => n14
                           );
   U16 : MUX2_X1 port map( A => Q_17_port, B => data(17), S => enable, Z => n15
                           );
   U17 : MUX2_X1 port map( A => Q_16_port, B => data(16), S => enable, Z => n16
                           );
   U18 : MUX2_X1 port map( A => Q_15_port, B => data(15), S => enable, Z => n17
                           );
   U19 : MUX2_X1 port map( A => Q_14_port, B => data(14), S => enable, Z => n18
                           );
   U20 : MUX2_X1 port map( A => Q_13_port, B => data(13), S => enable, Z => n19
                           );
   U21 : MUX2_X1 port map( A => Q_12_port, B => data(12), S => enable, Z => n20
                           );
   U22 : MUX2_X1 port map( A => Q_11_port, B => data(11), S => enable, Z => n21
                           );
   U23 : MUX2_X1 port map( A => Q_10_port, B => data(10), S => enable, Z => n22
                           );
   U24 : MUX2_X1 port map( A => Q_9_port, B => data(9), S => enable, Z => n23);
   U25 : MUX2_X1 port map( A => Q_8_port, B => data(8), S => enable, Z => n24);
   U26 : MUX2_X1 port map( A => Q_7_port, B => data(7), S => enable, Z => n25);
   U27 : MUX2_X1 port map( A => Q_6_port, B => data(6), S => enable, Z => n26);
   U28 : MUX2_X1 port map( A => Q_5_port, B => data(5), S => enable, Z => n27);
   U29 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n28);
   U30 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n29);
   U31 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n30);
   U32 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n31);
   U33 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n32);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N32_4 is

   port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end registro_N32_4;

architecture SYN_behaviour of registro_N32_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , net43347, net43348, net43349, net43350, net43351, net43352, net43353, 
      net43354, net43355, net43356, net43357, net43358, net43359, net43360, 
      net43361, net43362, net43363, net43364, net43365, net43366, net43367, 
      net43368, net43369, net43370, net43371, net43372, net43373, net43374, 
      net43375, net43376, net43377, net43378 : std_logic;

begin
   Q <= ( Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => clock, RN => clear, Q => 
                           Q_31_port, QN => net43378);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => clock, RN => clear, Q => 
                           Q_30_port, QN => net43377);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => clock, RN => clear, Q => 
                           Q_29_port, QN => net43376);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => clock, RN => clear, Q => 
                           Q_28_port, QN => net43375);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => clock, RN => clear, Q => 
                           Q_27_port, QN => net43374);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => clock, RN => clear, Q => 
                           Q_26_port, QN => net43373);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => clock, RN => clear, Q => 
                           Q_25_port, QN => net43372);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => clock, RN => clear, Q => 
                           Q_24_port, QN => net43371);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => clock, RN => clear, Q => 
                           Q_23_port, QN => net43370);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => clock, RN => clear, Q => 
                           Q_22_port, QN => net43369);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => clock, RN => clear, Q => 
                           Q_21_port, QN => net43368);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => clock, RN => clear, Q => 
                           Q_20_port, QN => net43367);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => clock, RN => clear, Q => 
                           Q_19_port, QN => net43366);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => clock, RN => clear, Q => 
                           Q_18_port, QN => net43365);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => clock, RN => clear, Q => 
                           Q_17_port, QN => net43364);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => clock, RN => clear, Q => 
                           Q_16_port, QN => net43363);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => clock, RN => clear, Q => 
                           Q_15_port, QN => net43362);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => clock, RN => clear, Q => 
                           Q_14_port, QN => net43361);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => clock, RN => clear, Q => 
                           Q_13_port, QN => net43360);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => clock, RN => clear, Q => 
                           Q_12_port, QN => net43359);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => clock, RN => clear, Q => 
                           Q_11_port, QN => net43358);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => clock, RN => clear, Q => 
                           Q_10_port, QN => net43357);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => clock, RN => clear, Q => 
                           Q_9_port, QN => net43356);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => clock, RN => clear, Q => 
                           Q_8_port, QN => net43355);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => clock, RN => clear, Q => 
                           Q_7_port, QN => net43354);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => clock, RN => clear, Q => 
                           Q_6_port, QN => net43353);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => clock, RN => clear, Q => 
                           Q_5_port, QN => net43352);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43351);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43350);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43349);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43348);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43347);
   U2 : MUX2_X1 port map( A => Q_31_port, B => data(31), S => enable, Z => n1);
   U3 : MUX2_X1 port map( A => Q_30_port, B => data(30), S => enable, Z => n2);
   U4 : MUX2_X1 port map( A => Q_29_port, B => data(29), S => enable, Z => n3);
   U5 : MUX2_X1 port map( A => Q_28_port, B => data(28), S => enable, Z => n4);
   U6 : MUX2_X1 port map( A => Q_27_port, B => data(27), S => enable, Z => n5);
   U7 : MUX2_X1 port map( A => Q_26_port, B => data(26), S => enable, Z => n6);
   U8 : MUX2_X1 port map( A => Q_25_port, B => data(25), S => enable, Z => n7);
   U9 : MUX2_X1 port map( A => Q_24_port, B => data(24), S => enable, Z => n8);
   U10 : MUX2_X1 port map( A => Q_23_port, B => data(23), S => enable, Z => n9)
                           ;
   U11 : MUX2_X1 port map( A => Q_22_port, B => data(22), S => enable, Z => n10
                           );
   U12 : MUX2_X1 port map( A => Q_21_port, B => data(21), S => enable, Z => n11
                           );
   U13 : MUX2_X1 port map( A => Q_20_port, B => data(20), S => enable, Z => n12
                           );
   U14 : MUX2_X1 port map( A => Q_19_port, B => data(19), S => enable, Z => n13
                           );
   U15 : MUX2_X1 port map( A => Q_18_port, B => data(18), S => enable, Z => n14
                           );
   U16 : MUX2_X1 port map( A => Q_17_port, B => data(17), S => enable, Z => n15
                           );
   U17 : MUX2_X1 port map( A => Q_16_port, B => data(16), S => enable, Z => n16
                           );
   U18 : MUX2_X1 port map( A => Q_15_port, B => data(15), S => enable, Z => n17
                           );
   U19 : MUX2_X1 port map( A => Q_14_port, B => data(14), S => enable, Z => n18
                           );
   U20 : MUX2_X1 port map( A => Q_13_port, B => data(13), S => enable, Z => n19
                           );
   U21 : MUX2_X1 port map( A => Q_12_port, B => data(12), S => enable, Z => n20
                           );
   U22 : MUX2_X1 port map( A => Q_11_port, B => data(11), S => enable, Z => n21
                           );
   U23 : MUX2_X1 port map( A => Q_10_port, B => data(10), S => enable, Z => n22
                           );
   U24 : MUX2_X1 port map( A => Q_9_port, B => data(9), S => enable, Z => n23);
   U25 : MUX2_X1 port map( A => Q_8_port, B => data(8), S => enable, Z => n24);
   U26 : MUX2_X1 port map( A => Q_7_port, B => data(7), S => enable, Z => n25);
   U27 : MUX2_X1 port map( A => Q_6_port, B => data(6), S => enable, Z => n26);
   U28 : MUX2_X1 port map( A => Q_5_port, B => data(5), S => enable, Z => n27);
   U29 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n28);
   U30 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n29);
   U31 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n30);
   U32 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n31);
   U33 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n32);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N32_3 is

   port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end registro_N32_3;

architecture SYN_behaviour of registro_N32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , net43315, net43316, net43317, net43318, net43319, net43320, net43321, 
      net43322, net43323, net43324, net43325, net43326, net43327, net43328, 
      net43329, net43330, net43331, net43332, net43333, net43334, net43335, 
      net43336, net43337, net43338, net43339, net43340, net43341, net43342, 
      net43343, net43344, net43345, net43346 : std_logic;

begin
   Q <= ( Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => clock, RN => clear, Q => 
                           Q_31_port, QN => net43346);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => clock, RN => clear, Q => 
                           Q_30_port, QN => net43345);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => clock, RN => clear, Q => 
                           Q_29_port, QN => net43344);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => clock, RN => clear, Q => 
                           Q_28_port, QN => net43343);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => clock, RN => clear, Q => 
                           Q_27_port, QN => net43342);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => clock, RN => clear, Q => 
                           Q_26_port, QN => net43341);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => clock, RN => clear, Q => 
                           Q_25_port, QN => net43340);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => clock, RN => clear, Q => 
                           Q_24_port, QN => net43339);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => clock, RN => clear, Q => 
                           Q_23_port, QN => net43338);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => clock, RN => clear, Q => 
                           Q_22_port, QN => net43337);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => clock, RN => clear, Q => 
                           Q_21_port, QN => net43336);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => clock, RN => clear, Q => 
                           Q_20_port, QN => net43335);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => clock, RN => clear, Q => 
                           Q_19_port, QN => net43334);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => clock, RN => clear, Q => 
                           Q_18_port, QN => net43333);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => clock, RN => clear, Q => 
                           Q_17_port, QN => net43332);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => clock, RN => clear, Q => 
                           Q_16_port, QN => net43331);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => clock, RN => clear, Q => 
                           Q_15_port, QN => net43330);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => clock, RN => clear, Q => 
                           Q_14_port, QN => net43329);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => clock, RN => clear, Q => 
                           Q_13_port, QN => net43328);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => clock, RN => clear, Q => 
                           Q_12_port, QN => net43327);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => clock, RN => clear, Q => 
                           Q_11_port, QN => net43326);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => clock, RN => clear, Q => 
                           Q_10_port, QN => net43325);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => clock, RN => clear, Q => 
                           Q_9_port, QN => net43324);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => clock, RN => clear, Q => 
                           Q_8_port, QN => net43323);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => clock, RN => clear, Q => 
                           Q_7_port, QN => net43322);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => clock, RN => clear, Q => 
                           Q_6_port, QN => net43321);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => clock, RN => clear, Q => 
                           Q_5_port, QN => net43320);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43319);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43318);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43317);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43316);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43315);
   U2 : MUX2_X1 port map( A => Q_31_port, B => data(31), S => enable, Z => n1);
   U3 : MUX2_X1 port map( A => Q_30_port, B => data(30), S => enable, Z => n2);
   U4 : MUX2_X1 port map( A => Q_29_port, B => data(29), S => enable, Z => n3);
   U5 : MUX2_X1 port map( A => Q_28_port, B => data(28), S => enable, Z => n4);
   U6 : MUX2_X1 port map( A => Q_27_port, B => data(27), S => enable, Z => n5);
   U7 : MUX2_X1 port map( A => Q_26_port, B => data(26), S => enable, Z => n6);
   U8 : MUX2_X1 port map( A => Q_25_port, B => data(25), S => enable, Z => n7);
   U9 : MUX2_X1 port map( A => Q_24_port, B => data(24), S => enable, Z => n8);
   U10 : MUX2_X1 port map( A => Q_23_port, B => data(23), S => enable, Z => n9)
                           ;
   U11 : MUX2_X1 port map( A => Q_22_port, B => data(22), S => enable, Z => n10
                           );
   U12 : MUX2_X1 port map( A => Q_21_port, B => data(21), S => enable, Z => n11
                           );
   U13 : MUX2_X1 port map( A => Q_20_port, B => data(20), S => enable, Z => n12
                           );
   U14 : MUX2_X1 port map( A => Q_19_port, B => data(19), S => enable, Z => n13
                           );
   U15 : MUX2_X1 port map( A => Q_18_port, B => data(18), S => enable, Z => n14
                           );
   U16 : MUX2_X1 port map( A => Q_17_port, B => data(17), S => enable, Z => n15
                           );
   U17 : MUX2_X1 port map( A => Q_16_port, B => data(16), S => enable, Z => n16
                           );
   U18 : MUX2_X1 port map( A => Q_15_port, B => data(15), S => enable, Z => n17
                           );
   U19 : MUX2_X1 port map( A => Q_14_port, B => data(14), S => enable, Z => n18
                           );
   U20 : MUX2_X1 port map( A => Q_13_port, B => data(13), S => enable, Z => n19
                           );
   U21 : MUX2_X1 port map( A => Q_12_port, B => data(12), S => enable, Z => n20
                           );
   U22 : MUX2_X1 port map( A => Q_11_port, B => data(11), S => enable, Z => n21
                           );
   U23 : MUX2_X1 port map( A => Q_10_port, B => data(10), S => enable, Z => n22
                           );
   U24 : MUX2_X1 port map( A => Q_9_port, B => data(9), S => enable, Z => n23);
   U25 : MUX2_X1 port map( A => Q_8_port, B => data(8), S => enable, Z => n24);
   U26 : MUX2_X1 port map( A => Q_7_port, B => data(7), S => enable, Z => n25);
   U27 : MUX2_X1 port map( A => Q_6_port, B => data(6), S => enable, Z => n26);
   U28 : MUX2_X1 port map( A => Q_5_port, B => data(5), S => enable, Z => n27);
   U29 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n28);
   U30 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n29);
   U31 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n30);
   U32 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n31);
   U33 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n32);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N32_2 is

   port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end registro_N32_2;

architecture SYN_behaviour of registro_N32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , net43283, net43284, net43285, net43286, net43287, net43288, net43289, 
      net43290, net43291, net43292, net43293, net43294, net43295, net43296, 
      net43297, net43298, net43299, net43300, net43301, net43302, net43303, 
      net43304, net43305, net43306, net43307, net43308, net43309, net43310, 
      net43311, net43312, net43313, net43314 : std_logic;

begin
   Q <= ( Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => clock, RN => clear, Q => 
                           Q_31_port, QN => net43314);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => clock, RN => clear, Q => 
                           Q_30_port, QN => net43313);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => clock, RN => clear, Q => 
                           Q_29_port, QN => net43312);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => clock, RN => clear, Q => 
                           Q_28_port, QN => net43311);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => clock, RN => clear, Q => 
                           Q_27_port, QN => net43310);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => clock, RN => clear, Q => 
                           Q_26_port, QN => net43309);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => clock, RN => clear, Q => 
                           Q_25_port, QN => net43308);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => clock, RN => clear, Q => 
                           Q_24_port, QN => net43307);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => clock, RN => clear, Q => 
                           Q_23_port, QN => net43306);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => clock, RN => clear, Q => 
                           Q_22_port, QN => net43305);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => clock, RN => clear, Q => 
                           Q_21_port, QN => net43304);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => clock, RN => clear, Q => 
                           Q_20_port, QN => net43303);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => clock, RN => clear, Q => 
                           Q_19_port, QN => net43302);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => clock, RN => clear, Q => 
                           Q_18_port, QN => net43301);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => clock, RN => clear, Q => 
                           Q_17_port, QN => net43300);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => clock, RN => clear, Q => 
                           Q_16_port, QN => net43299);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => clock, RN => clear, Q => 
                           Q_15_port, QN => net43298);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => clock, RN => clear, Q => 
                           Q_14_port, QN => net43297);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => clock, RN => clear, Q => 
                           Q_13_port, QN => net43296);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => clock, RN => clear, Q => 
                           Q_12_port, QN => net43295);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => clock, RN => clear, Q => 
                           Q_11_port, QN => net43294);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => clock, RN => clear, Q => 
                           Q_10_port, QN => net43293);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => clock, RN => clear, Q => 
                           Q_9_port, QN => net43292);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => clock, RN => clear, Q => 
                           Q_8_port, QN => net43291);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => clock, RN => clear, Q => 
                           Q_7_port, QN => net43290);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => clock, RN => clear, Q => 
                           Q_6_port, QN => net43289);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => clock, RN => clear, Q => 
                           Q_5_port, QN => net43288);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43287);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43286);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43285);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43284);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43283);
   U2 : MUX2_X1 port map( A => Q_31_port, B => data(31), S => enable, Z => n1);
   U3 : MUX2_X1 port map( A => Q_30_port, B => data(30), S => enable, Z => n2);
   U4 : MUX2_X1 port map( A => Q_29_port, B => data(29), S => enable, Z => n3);
   U5 : MUX2_X1 port map( A => Q_28_port, B => data(28), S => enable, Z => n4);
   U6 : MUX2_X1 port map( A => Q_27_port, B => data(27), S => enable, Z => n5);
   U7 : MUX2_X1 port map( A => Q_26_port, B => data(26), S => enable, Z => n6);
   U8 : MUX2_X1 port map( A => Q_25_port, B => data(25), S => enable, Z => n7);
   U9 : MUX2_X1 port map( A => Q_24_port, B => data(24), S => enable, Z => n8);
   U10 : MUX2_X1 port map( A => Q_23_port, B => data(23), S => enable, Z => n9)
                           ;
   U11 : MUX2_X1 port map( A => Q_22_port, B => data(22), S => enable, Z => n10
                           );
   U12 : MUX2_X1 port map( A => Q_21_port, B => data(21), S => enable, Z => n11
                           );
   U13 : MUX2_X1 port map( A => Q_20_port, B => data(20), S => enable, Z => n12
                           );
   U14 : MUX2_X1 port map( A => Q_19_port, B => data(19), S => enable, Z => n13
                           );
   U15 : MUX2_X1 port map( A => Q_18_port, B => data(18), S => enable, Z => n14
                           );
   U16 : MUX2_X1 port map( A => Q_17_port, B => data(17), S => enable, Z => n15
                           );
   U17 : MUX2_X1 port map( A => Q_16_port, B => data(16), S => enable, Z => n16
                           );
   U18 : MUX2_X1 port map( A => Q_15_port, B => data(15), S => enable, Z => n17
                           );
   U19 : MUX2_X1 port map( A => Q_14_port, B => data(14), S => enable, Z => n18
                           );
   U20 : MUX2_X1 port map( A => Q_13_port, B => data(13), S => enable, Z => n19
                           );
   U21 : MUX2_X1 port map( A => Q_12_port, B => data(12), S => enable, Z => n20
                           );
   U22 : MUX2_X1 port map( A => Q_11_port, B => data(11), S => enable, Z => n21
                           );
   U23 : MUX2_X1 port map( A => Q_10_port, B => data(10), S => enable, Z => n22
                           );
   U24 : MUX2_X1 port map( A => Q_9_port, B => data(9), S => enable, Z => n23);
   U25 : MUX2_X1 port map( A => Q_8_port, B => data(8), S => enable, Z => n24);
   U26 : MUX2_X1 port map( A => Q_7_port, B => data(7), S => enable, Z => n25);
   U27 : MUX2_X1 port map( A => Q_6_port, B => data(6), S => enable, Z => n26);
   U28 : MUX2_X1 port map( A => Q_5_port, B => data(5), S => enable, Z => n27);
   U29 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n28);
   U30 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n29);
   U31 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n30);
   U32 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n31);
   U33 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n32);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N32_1 is

   port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end registro_N32_1;

architecture SYN_behaviour of registro_N32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n1,
      n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, 
      n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32
      , net43251, net43252, net43253, net43254, net43255, net43256, net43257, 
      net43258, net43259, net43260, net43261, net43262, net43263, net43264, 
      net43265, net43266, net43267, net43268, net43269, net43270, net43271, 
      net43272, net43273, net43274, net43275, net43276, net43277, net43278, 
      net43279, net43280, net43281, net43282 : std_logic;

begin
   Q <= ( Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_31_inst : DFFR_X1 port map( D => n1, CK => clock, RN => clear, Q => 
                           Q_31_port, QN => net43282);
   Q_reg_30_inst : DFFR_X1 port map( D => n2, CK => clock, RN => clear, Q => 
                           Q_30_port, QN => net43281);
   Q_reg_29_inst : DFFR_X1 port map( D => n3, CK => clock, RN => clear, Q => 
                           Q_29_port, QN => net43280);
   Q_reg_28_inst : DFFR_X1 port map( D => n4, CK => clock, RN => clear, Q => 
                           Q_28_port, QN => net43279);
   Q_reg_27_inst : DFFR_X1 port map( D => n5, CK => clock, RN => clear, Q => 
                           Q_27_port, QN => net43278);
   Q_reg_26_inst : DFFR_X1 port map( D => n6, CK => clock, RN => clear, Q => 
                           Q_26_port, QN => net43277);
   Q_reg_25_inst : DFFR_X1 port map( D => n7, CK => clock, RN => clear, Q => 
                           Q_25_port, QN => net43276);
   Q_reg_24_inst : DFFR_X1 port map( D => n8, CK => clock, RN => clear, Q => 
                           Q_24_port, QN => net43275);
   Q_reg_23_inst : DFFR_X1 port map( D => n9, CK => clock, RN => clear, Q => 
                           Q_23_port, QN => net43274);
   Q_reg_22_inst : DFFR_X1 port map( D => n10, CK => clock, RN => clear, Q => 
                           Q_22_port, QN => net43273);
   Q_reg_21_inst : DFFR_X1 port map( D => n11, CK => clock, RN => clear, Q => 
                           Q_21_port, QN => net43272);
   Q_reg_20_inst : DFFR_X1 port map( D => n12, CK => clock, RN => clear, Q => 
                           Q_20_port, QN => net43271);
   Q_reg_19_inst : DFFR_X1 port map( D => n13, CK => clock, RN => clear, Q => 
                           Q_19_port, QN => net43270);
   Q_reg_18_inst : DFFR_X1 port map( D => n14, CK => clock, RN => clear, Q => 
                           Q_18_port, QN => net43269);
   Q_reg_17_inst : DFFR_X1 port map( D => n15, CK => clock, RN => clear, Q => 
                           Q_17_port, QN => net43268);
   Q_reg_16_inst : DFFR_X1 port map( D => n16, CK => clock, RN => clear, Q => 
                           Q_16_port, QN => net43267);
   Q_reg_15_inst : DFFR_X1 port map( D => n17, CK => clock, RN => clear, Q => 
                           Q_15_port, QN => net43266);
   Q_reg_14_inst : DFFR_X1 port map( D => n18, CK => clock, RN => clear, Q => 
                           Q_14_port, QN => net43265);
   Q_reg_13_inst : DFFR_X1 port map( D => n19, CK => clock, RN => clear, Q => 
                           Q_13_port, QN => net43264);
   Q_reg_12_inst : DFFR_X1 port map( D => n20, CK => clock, RN => clear, Q => 
                           Q_12_port, QN => net43263);
   Q_reg_11_inst : DFFR_X1 port map( D => n21, CK => clock, RN => clear, Q => 
                           Q_11_port, QN => net43262);
   Q_reg_10_inst : DFFR_X1 port map( D => n22, CK => clock, RN => clear, Q => 
                           Q_10_port, QN => net43261);
   Q_reg_9_inst : DFFR_X1 port map( D => n23, CK => clock, RN => clear, Q => 
                           Q_9_port, QN => net43260);
   Q_reg_8_inst : DFFR_X1 port map( D => n24, CK => clock, RN => clear, Q => 
                           Q_8_port, QN => net43259);
   Q_reg_7_inst : DFFR_X1 port map( D => n25, CK => clock, RN => clear, Q => 
                           Q_7_port, QN => net43258);
   Q_reg_6_inst : DFFR_X1 port map( D => n26, CK => clock, RN => clear, Q => 
                           Q_6_port, QN => net43257);
   Q_reg_5_inst : DFFR_X1 port map( D => n27, CK => clock, RN => clear, Q => 
                           Q_5_port, QN => net43256);
   Q_reg_4_inst : DFFR_X1 port map( D => n28, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43255);
   Q_reg_3_inst : DFFR_X1 port map( D => n29, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43254);
   Q_reg_2_inst : DFFR_X1 port map( D => n30, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43253);
   Q_reg_1_inst : DFFR_X1 port map( D => n31, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43252);
   Q_reg_0_inst : DFFR_X1 port map( D => n32, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43251);
   U2 : MUX2_X1 port map( A => Q_31_port, B => data(31), S => enable, Z => n1);
   U3 : MUX2_X1 port map( A => Q_30_port, B => data(30), S => enable, Z => n2);
   U4 : MUX2_X1 port map( A => Q_29_port, B => data(29), S => enable, Z => n3);
   U5 : MUX2_X1 port map( A => Q_28_port, B => data(28), S => enable, Z => n4);
   U6 : MUX2_X1 port map( A => Q_27_port, B => data(27), S => enable, Z => n5);
   U7 : MUX2_X1 port map( A => Q_26_port, B => data(26), S => enable, Z => n6);
   U8 : MUX2_X1 port map( A => Q_25_port, B => data(25), S => enable, Z => n7);
   U9 : MUX2_X1 port map( A => Q_24_port, B => data(24), S => enable, Z => n8);
   U10 : MUX2_X1 port map( A => Q_23_port, B => data(23), S => enable, Z => n9)
                           ;
   U11 : MUX2_X1 port map( A => Q_22_port, B => data(22), S => enable, Z => n10
                           );
   U12 : MUX2_X1 port map( A => Q_21_port, B => data(21), S => enable, Z => n11
                           );
   U13 : MUX2_X1 port map( A => Q_20_port, B => data(20), S => enable, Z => n12
                           );
   U14 : MUX2_X1 port map( A => Q_19_port, B => data(19), S => enable, Z => n13
                           );
   U15 : MUX2_X1 port map( A => Q_18_port, B => data(18), S => enable, Z => n14
                           );
   U16 : MUX2_X1 port map( A => Q_17_port, B => data(17), S => enable, Z => n15
                           );
   U17 : MUX2_X1 port map( A => Q_16_port, B => data(16), S => enable, Z => n16
                           );
   U18 : MUX2_X1 port map( A => Q_15_port, B => data(15), S => enable, Z => n17
                           );
   U19 : MUX2_X1 port map( A => Q_14_port, B => data(14), S => enable, Z => n18
                           );
   U20 : MUX2_X1 port map( A => Q_13_port, B => data(13), S => enable, Z => n19
                           );
   U21 : MUX2_X1 port map( A => Q_12_port, B => data(12), S => enable, Z => n20
                           );
   U22 : MUX2_X1 port map( A => Q_11_port, B => data(11), S => enable, Z => n21
                           );
   U23 : MUX2_X1 port map( A => Q_10_port, B => data(10), S => enable, Z => n22
                           );
   U24 : MUX2_X1 port map( A => Q_9_port, B => data(9), S => enable, Z => n23);
   U25 : MUX2_X1 port map( A => Q_8_port, B => data(8), S => enable, Z => n24);
   U26 : MUX2_X1 port map( A => Q_7_port, B => data(7), S => enable, Z => n25);
   U27 : MUX2_X1 port map( A => Q_6_port, B => data(6), S => enable, Z => n26);
   U28 : MUX2_X1 port map( A => Q_5_port, B => data(5), S => enable, Z => n27);
   U29 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n28);
   U30 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n29);
   U31 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n30);
   U32 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n31);
   U33 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n32);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_N32_4 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end mux21_N32_4;

architecture SYN_behavioural of mux21_N32_4 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component MUX2_X2
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X2 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U2 : MUX2_X2 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U3 : MUX2_X2 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U4 : MUX2_X2 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U5 : MUX2_X2 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U6 : MUX2_X2 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U7 : MUX2_X2 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U8 : MUX2_X2 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U9 : MUX2_X2 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U10 : MUX2_X2 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U11 : MUX2_X2 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U12 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U13 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U14 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U15 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U16 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U17 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U18 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U19 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U20 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U21 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U22 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U23 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U24 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U25 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U26 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U27 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U28 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U29 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U30 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U31 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_N32_3 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end mux21_N32_3;

architecture SYN_behavioural of mux21_N32_3 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n9, n10, n11, n12, n1, n3, n5, n7 : std_logic;

begin
   
   U1 : INV_X1 port map( A => n10, ZN => n1);
   U2 : INV_X8 port map( A => n1, ZN => Y(2));
   U3 : INV_X1 port map( A => n9, ZN => n3);
   U4 : INV_X8 port map( A => n3, ZN => Y(3));
   U5 : INV_X1 port map( A => n12, ZN => n5);
   U6 : INV_X8 port map( A => n5, ZN => Y(0));
   U7 : INV_X1 port map( A => n11, ZN => n7);
   U8 : INV_X8 port map( A => n7, ZN => Y(1));
   U9 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U10 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U11 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U12 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U13 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U14 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U15 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => n9);
   U16 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U17 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U18 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => n10);
   U19 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U20 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U21 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U22 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U23 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U24 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U25 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U26 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U27 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U28 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U29 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => n11);
   U30 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U31 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U32 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U33 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U34 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U35 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U36 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U37 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U38 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U39 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U40 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => n12);

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_N32_2 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end mux21_N32_2;

architecture SYN_behavioural of mux21_N32_2 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U2 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U3 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U4 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U5 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U6 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U7 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U8 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U9 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U10 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U11 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U12 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U13 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U14 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U15 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U16 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U17 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U18 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U19 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U20 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U21 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U22 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U23 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U26 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U27 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U28 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U29 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U30 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U31 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_N32_1 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end mux21_N32_1;

architecture SYN_behavioural of mux21_N32_1 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U2 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U3 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U4 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U5 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U6 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U7 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U8 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U9 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U10 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U11 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U12 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U13 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U14 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U15 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U16 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U17 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U18 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U19 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U20 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U21 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U22 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U23 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U26 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U27 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U28 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U29 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U30 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U31 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_generic_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (3 downto 0));

end mux21_generic_NBIT4_0;

architecture SYN_behavioural of mux21_generic_NBIT4_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => B(3), B => A(3), S => SEL, Z => Y(3));
   U2 : MUX2_X1 port map( A => B(2), B => A(2), S => SEL, Z => Y(2));
   U3 : MUX2_X1 port map( A => B(1), B => A(1), S => SEL, Z => Y(1));
   U4 : MUX2_X1 port map( A => B(0), B => A(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : out 
         std_logic_vector (3 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT4_0;

architecture SYN_structural of RCA_GEN_NBIT4_0 is

   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_64
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_3_port, CTMP_2_port, CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_64 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_63 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_62 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_61 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PGnet_0 is

   port( A, B, C : in std_logic;  P, G : out std_logic);

end PGnet_0;

architecture SYN_beh of PGnet_0 is

   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : XOR2_X1 port map( A => B, B => A, Z => P);
   U2 : AND2_X1 port map( A1 => B, A2 => A, ZN => G);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity carry_select_N4_0 is

   port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : out
         std_logic_vector (3 downto 0));

end carry_select_N4_0;

architecture SYN_beh of carry_select_N4_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component mux21_generic_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component RCA_GEN_NBIT4_15
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   component RCA_GEN_NBIT4_0
      port( A, B : in std_logic_vector (3 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (3 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, sel, S0_3_port, S0_2_port, S0_1_port, 
      S0_0_port, S1_3_port, S1_2_port, S1_1_port, S1_0_port, net2289, net2290 :
      std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   RCA1 : RCA_GEN_NBIT4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic0_port, S(3) => 
                           S0_3_port, S(2) => S0_2_port, S(1) => S0_1_port, 
                           S(0) => S0_0_port, Co => net2290);
   RCA2 : RCA_GEN_NBIT4_15 port map( A(3) => A(3), A(2) => A(2), A(1) => A(1), 
                           A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1) => 
                           B(1), B(0) => B(0), Ci => X_Logic1_port, S(3) => 
                           S1_3_port, S(2) => S1_2_port, S(1) => S1_1_port, 
                           S(0) => S1_0_port, Co => net2289);
   MUX1 : mux21_generic_NBIT4_0 port map( A(3) => S0_3_port, A(2) => S0_2_port,
                           A(1) => S0_1_port, A(0) => S0_0_port, B(3) => 
                           S1_3_port, B(2) => S1_2_port, B(1) => S1_1_port, 
                           B(0) => S1_0_port, SEL => sel, Y(3) => S(3), Y(2) =>
                           S(2), Y(1) => S(1), Y(0) => S(0));
   U3 : INV_X1 port map( A => Cin, ZN => sel);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity PG_0 is

   port( A, B, C, D : in std_logic;  P, G : out std_logic);

end PG_0;

architecture SYN_beh of PG_0 is

   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1 : std_logic;

begin
   
   U1 : AND2_X1 port map( A1 => B, A2 => A, ZN => P);
   U2 : INV_X1 port map( A => n1, ZN => G);
   U3 : AOI21_X1 port map( B1 => D, B2 => A, A => C, ZN => n1);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sparse_tree_carry_gen_4bits_0 is

   port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, G :
         out std_logic);

end sparse_tree_carry_gen_4bits_0;

architecture SYN_beh of sparse_tree_carry_gen_4bits_0 is

   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component PG_22
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_23
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_24
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_22
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_23
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   component PGnet_0
      port( A, B, C : in std_logic;  P, G : out std_logic);
   end component;
   
   signal X_Logic0_port, P0_3_port, P0_2_port, P0_1_port, P0_0_port, G0_3_port,
      G0_2_port, G0_1_port, G0_0_port, G1_1_port, G1_0_port, P1_1_port, 
      P1_0_port, n1, n2, n3 : std_logic;

begin
   
   X_Logic0_port <= '0';
   pg1_1 : PGnet_0 port map( A => A(1), B => B(1), C => X_Logic0_port, P => 
                           P0_1_port, G => G0_1_port);
   pg1_2 : PGnet_23 port map( A => A(2), B => B(2), C => X_Logic0_port, P => 
                           P0_2_port, G => G0_2_port);
   pg1_3 : PGnet_22 port map( A => A(3), B => B(3), C => X_Logic0_port, P => 
                           P0_3_port, G => G0_3_port);
   pg2_0 : PG_24 port map( A => P0_1_port, B => P0_0_port, C => G0_1_port, D =>
                           G0_0_port, P => P1_0_port, G => G1_0_port);
   pg2_1 : PG_23 port map( A => P0_3_port, B => P0_2_port, C => G0_3_port, D =>
                           G0_2_port, P => P1_1_port, G => G1_1_port);
   pgg : PG_22 port map( A => P1_1_port, B => P1_0_port, C => G1_1_port, D => 
                           G1_0_port, P => P, G => G);
   U2 : XOR2_X1 port map( A => B(0), B => A(0), Z => P0_0_port);
   U3 : INV_X1 port map( A => n1, ZN => G0_0_port);
   U4 : AOI21_X1 port map( B1 => B(0), B2 => A(0), A => n2, ZN => n1);
   U5 : INV_X1 port map( A => n3, ZN => n2);
   U6 : OAI21_X1 port map( B1 => A(0), B2 => B(0), A => c_in, ZN => n3);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sum_generator_N32_N_carry4 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector (8
         downto 0);  Sum : out std_logic_vector (31 downto 0));

end sum_generator_N32_N_carry4;

architecture SYN_behaviour of sum_generator_N32_N_carry4 is

   component carry_select_N4_1
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_2
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_3
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_4
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_5
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_6
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_7
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;
   
   component carry_select_N4_0
      port( A, B : in std_logic_vector (3 downto 0);  Cin : in std_logic;  S : 
            out std_logic_vector (3 downto 0));
   end component;

begin
   
   CBLOCk_0 : carry_select_N4_0 port map( A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(3) => B(3), B(2) => B(2), B(1)
                           => B(1), B(0) => B(0), Cin => Ci(0), S(3) => Sum(3),
                           S(2) => Sum(2), S(1) => Sum(1), S(0) => Sum(0));
   CBLOCk_1 : carry_select_N4_7 port map( A(3) => A(7), A(2) => A(6), A(1) => 
                           A(5), A(0) => A(4), B(3) => B(7), B(2) => B(6), B(1)
                           => B(5), B(0) => B(4), Cin => Ci(1), S(3) => Sum(7),
                           S(2) => Sum(6), S(1) => Sum(5), S(0) => Sum(4));
   CBLOCk_2 : carry_select_N4_6 port map( A(3) => A(11), A(2) => A(10), A(1) =>
                           A(9), A(0) => A(8), B(3) => B(11), B(2) => B(10), 
                           B(1) => B(9), B(0) => B(8), Cin => Ci(2), S(3) => 
                           Sum(11), S(2) => Sum(10), S(1) => Sum(9), S(0) => 
                           Sum(8));
   CBLOCk_3 : carry_select_N4_5 port map( A(3) => A(15), A(2) => A(14), A(1) =>
                           A(13), A(0) => A(12), B(3) => B(15), B(2) => B(14), 
                           B(1) => B(13), B(0) => B(12), Cin => Ci(3), S(3) => 
                           Sum(15), S(2) => Sum(14), S(1) => Sum(13), S(0) => 
                           Sum(12));
   CBLOCk_4 : carry_select_N4_4 port map( A(3) => A(19), A(2) => A(18), A(1) =>
                           A(17), A(0) => A(16), B(3) => B(19), B(2) => B(18), 
                           B(1) => B(17), B(0) => B(16), Cin => Ci(4), S(3) => 
                           Sum(19), S(2) => Sum(18), S(1) => Sum(17), S(0) => 
                           Sum(16));
   CBLOCk_5 : carry_select_N4_3 port map( A(3) => A(23), A(2) => A(22), A(1) =>
                           A(21), A(0) => A(20), B(3) => B(23), B(2) => B(22), 
                           B(1) => B(21), B(0) => B(20), Cin => Ci(5), S(3) => 
                           Sum(23), S(2) => Sum(22), S(1) => Sum(21), S(0) => 
                           Sum(20));
   CBLOCk_6 : carry_select_N4_2 port map( A(3) => A(27), A(2) => A(26), A(1) =>
                           A(25), A(0) => A(24), B(3) => B(27), B(2) => B(26), 
                           B(1) => B(25), B(0) => B(24), Cin => Ci(6), S(3) => 
                           Sum(27), S(2) => Sum(26), S(1) => Sum(25), S(0) => 
                           Sum(24));
   CBLOCk_7 : carry_select_N4_1 port map( A(3) => A(31), A(2) => A(30), A(1) =>
                           A(29), A(0) => A(28), B(3) => B(31), B(2) => B(30), 
                           B(1) => B(29), B(0) => B(28), Cin => Ci(7), S(3) => 
                           Sum(31), S(2) => Sum(30), S(1) => Sum(29), S(0) => 
                           Sum(28));

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity sparse_tree_carry_gen_N5 is

   port( A, B : in std_logic_vector (31 downto 0);  C0 : in std_logic;  Cout : 
         out std_logic_vector (7 downto 0));

end sparse_tree_carry_gen_N5;

architecture SYN_beh of sparse_tree_carry_gen_N5 is

   component PG_25
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_26
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_27
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_28
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_29
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_30
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_31
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_32
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_33
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_34
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_35
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_36
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_37
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_38
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_39
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_40
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_41
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_42
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_43
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component PG_0
      port( A, B, C, D : in std_logic;  P, G : out std_logic);
   end component;
   
   component sparse_tree_carry_gen_4bits_1
      port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, 
            G : out std_logic);
   end component;
   
   component sparse_tree_carry_gen_4bits_2
      port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, 
            G : out std_logic);
   end component;
   
   component sparse_tree_carry_gen_4bits_3
      port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, 
            G : out std_logic);
   end component;
   
   component sparse_tree_carry_gen_4bits_4
      port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, 
            G : out std_logic);
   end component;
   
   component sparse_tree_carry_gen_4bits_5
      port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, 
            G : out std_logic);
   end component;
   
   component sparse_tree_carry_gen_4bits_6
      port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, 
            G : out std_logic);
   end component;
   
   component sparse_tree_carry_gen_4bits_7
      port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, 
            G : out std_logic);
   end component;
   
   component sparse_tree_carry_gen_4bits_0
      port( A, B : in std_logic_vector (3 downto 0);  c_in : in std_logic;  P, 
            G : out std_logic);
   end component;
   
   signal Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, Cout_3_port, 
      Cout_2_port, Cout_1_port, Cout_0_port, G_2_7_port, G_2_6_port, G_1_7_port
      , G_1_5_port, G_1_3_port, G_0_7_port, G_0_6_port, G_0_5_port, G_0_4_port,
      G_0_3_port, G_0_2_port, G_0_1_port, P_2_7_port, P_2_6_port, P_2_3_port, 
      P_2_2_port, P_1_7_port, P_1_5_port, P_1_3_port, P_1_1_port, P_1_0_port, 
      P_0_7_port, P_0_6_port, P_0_5_port, P_0_4_port, P_0_3_port, P_0_2_port, 
      P_0_1_port, net2281, net2282, net2283, net2284, net2285, net2286, net2287
      , net2288 : std_logic;

begin
   Cout <= ( Cout_7_port, Cout_6_port, Cout_5_port, Cout_4_port, Cout_3_port, 
      Cout_2_port, Cout_1_port, Cout_0_port );
   
   pg4_0_0 : sparse_tree_carry_gen_4bits_0 port map( A(3) => A(3), A(2) => A(2)
                           , A(1) => A(1), A(0) => A(0), B(3) => B(3), B(2) => 
                           B(2), B(1) => B(1), B(0) => B(0), c_in => C0, P => 
                           P_1_0_port, G => Cout_0_port);
   pg4_0_1 : sparse_tree_carry_gen_4bits_7 port map( A(3) => A(7), A(2) => A(6)
                           , A(1) => A(5), A(0) => A(4), B(3) => B(7), B(2) => 
                           B(6), B(1) => B(5), B(0) => B(4), c_in => C0, P => 
                           P_0_1_port, G => G_0_1_port);
   pg4_0_2 : sparse_tree_carry_gen_4bits_6 port map( A(3) => A(11), A(2) => 
                           A(10), A(1) => A(9), A(0) => A(8), B(3) => B(11), 
                           B(2) => B(10), B(1) => B(9), B(0) => B(8), c_in => 
                           C0, P => P_0_2_port, G => G_0_2_port);
   pg4_0_3 : sparse_tree_carry_gen_4bits_5 port map( A(3) => A(15), A(2) => 
                           A(14), A(1) => A(13), A(0) => A(12), B(3) => B(15), 
                           B(2) => B(14), B(1) => B(13), B(0) => B(12), c_in =>
                           C0, P => P_0_3_port, G => G_0_3_port);
   pg4_0_4 : sparse_tree_carry_gen_4bits_4 port map( A(3) => A(19), A(2) => 
                           A(18), A(1) => A(17), A(0) => A(16), B(3) => B(19), 
                           B(2) => B(18), B(1) => B(17), B(0) => B(16), c_in =>
                           C0, P => P_0_4_port, G => G_0_4_port);
   pg4_0_5 : sparse_tree_carry_gen_4bits_3 port map( A(3) => A(23), A(2) => 
                           A(22), A(1) => A(21), A(0) => A(20), B(3) => B(23), 
                           B(2) => B(22), B(1) => B(21), B(0) => B(20), c_in =>
                           C0, P => P_0_5_port, G => G_0_5_port);
   pg4_0_6 : sparse_tree_carry_gen_4bits_2 port map( A(3) => A(27), A(2) => 
                           A(26), A(1) => A(25), A(0) => A(24), B(3) => B(27), 
                           B(2) => B(26), B(1) => B(25), B(0) => B(24), c_in =>
                           C0, P => P_0_6_port, G => G_0_6_port);
   pg4_0_7 : sparse_tree_carry_gen_4bits_1 port map( A(3) => A(31), A(2) => 
                           A(30), A(1) => A(29), A(0) => A(28), B(3) => B(31), 
                           B(2) => B(30), B(1) => B(29), B(0) => B(28), c_in =>
                           C0, P => P_0_7_port, G => G_0_7_port);
   pg1_1_0 : PG_0 port map( A => P_0_1_port, B => P_1_0_port, C => G_0_1_port, 
                           D => Cout_0_port, P => P_1_1_port, G => Cout_1_port)
                           ;
   pg1_1_1 : PG_43 port map( A => P_0_3_port, B => P_0_2_port, C => G_0_3_port,
                           D => G_0_2_port, P => P_1_3_port, G => G_1_3_port);
   pg1_1_2 : PG_42 port map( A => P_0_5_port, B => P_0_4_port, C => G_0_5_port,
                           D => G_0_4_port, P => P_1_5_port, G => G_1_5_port);
   pg1_1_3 : PG_41 port map( A => P_0_7_port, B => P_0_6_port, C => G_0_7_port,
                           D => G_0_6_port, P => P_1_7_port, G => G_1_7_port);
   gen2_2_0_2_1 : PG_40 port map( A => P_0_2_port, B => P_1_1_port, C => 
                           G_0_2_port, D => Cout_1_port, P => P_2_2_port, G => 
                           Cout_2_port);
   gen2_2_0_2_2 : PG_39 port map( A => P_0_2_port, B => P_1_0_port, C => 
                           G_0_2_port, D => Cout_0_port, P => P_2_2_port, G => 
                           Cout_2_port);
   gen2_2_0_3_1 : PG_38 port map( A => P_1_3_port, B => P_0_2_port, C => 
                           G_1_3_port, D => G_0_2_port, P => P_2_3_port, G => 
                           Cout_3_port);
   gen2_2_0_3_2 : PG_37 port map( A => P_1_3_port, B => P_1_1_port, C => 
                           G_1_3_port, D => Cout_1_port, P => P_2_3_port, G => 
                           Cout_3_port);
   gen2_2_1_6_1 : PG_36 port map( A => P_0_6_port, B => P_1_5_port, C => 
                           G_0_6_port, D => G_1_5_port, P => P_2_6_port, G => 
                           G_2_6_port);
   gen2_2_1_6_2 : PG_35 port map( A => P_0_6_port, B => P_0_4_port, C => 
                           G_0_6_port, D => G_0_4_port, P => P_2_6_port, G => 
                           G_2_6_port);
   gen2_2_1_7_1 : PG_34 port map( A => P_1_7_port, B => P_0_6_port, C => 
                           G_1_7_port, D => G_0_6_port, P => P_2_7_port, G => 
                           G_2_7_port);
   gen2_2_1_7_2 : PG_33 port map( A => P_1_7_port, B => P_1_5_port, C => 
                           G_1_7_port, D => G_1_5_port, P => P_2_7_port, G => 
                           G_2_7_port);
   gen2_3_0_4_1 : PG_32 port map( A => P_0_4_port, B => P_2_3_port, C => 
                           G_0_4_port, D => Cout_3_port, P => net2288, G => 
                           Cout_4_port);
   gen2_3_0_4_2 : PG_31 port map( A => P_0_4_port, B => P_2_2_port, C => 
                           G_0_4_port, D => Cout_2_port, P => net2287, G => 
                           Cout_4_port);
   gen2_3_0_5_1 : PG_30 port map( A => P_1_5_port, B => P_0_4_port, C => 
                           G_1_5_port, D => G_0_4_port, P => net2286, G => 
                           Cout_5_port);
   gen2_3_0_5_2 : PG_29 port map( A => P_1_5_port, B => P_2_3_port, C => 
                           G_1_5_port, D => Cout_3_port, P => net2285, G => 
                           Cout_5_port);
   gen2_3_0_6_1 : PG_28 port map( A => P_2_6_port, B => P_1_5_port, C => 
                           G_2_6_port, D => G_1_5_port, P => net2284, G => 
                           Cout_6_port);
   gen2_3_0_6_2 : PG_27 port map( A => P_2_6_port, B => P_0_4_port, C => 
                           G_2_6_port, D => G_0_4_port, P => net2283, G => 
                           Cout_6_port);
   gen2_3_0_7_1 : PG_26 port map( A => P_2_7_port, B => P_2_6_port, C => 
                           G_2_7_port, D => G_2_6_port, P => net2282, G => 
                           Cout_7_port);
   gen2_3_0_7_2 : PG_25 port map( A => P_2_7_port, B => P_1_5_port, C => 
                           G_2_7_port, D => G_1_5_port, P => net2281, G => 
                           Cout_7_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_6to1_n32 is

   port( A, B, C, D, E, F : in std_logic_vector (31 downto 0);  S : in 
         std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto 0)
         );

end MUX_6to1_n32;

architecture SYN_BEH of MUX_6to1_n32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74
      , n75, n76, n77, n78, n79, n80 : std_logic;

begin
   
   U1 : CLKBUF_X2 port map( A => n14, Z => n1);
   U2 : OR3_X1 port map( A1 => S(0), A2 => S(2), A3 => n79, ZN => n2);
   U3 : INV_X2 port map( A => n2, ZN => n3);
   U4 : OR3_X1 port map( A1 => n78, A2 => S(1), A3 => n80, ZN => n4);
   U5 : INV_X2 port map( A => n4, ZN => n5);
   U6 : OR3_X1 port map( A1 => S(1), A2 => S(2), A3 => n78, ZN => n6);
   U7 : INV_X2 port map( A => n6, ZN => n7);
   U8 : OR3_X1 port map( A1 => n78, A2 => S(2), A3 => n79, ZN => n8);
   U9 : INV_X2 port map( A => n8, ZN => n9);
   U10 : OR3_X1 port map( A1 => S(0), A2 => S(1), A3 => n80, ZN => n10);
   U11 : INV_X2 port map( A => n10, ZN => n11);
   U12 : NAND2_X1 port map( A1 => n12, A2 => n13, ZN => Y(9));
   U13 : AOI222_X1 port map( A1 => E(9), A2 => n11, B1 => A(9), B2 => n1, C1 =>
                           D(9), C2 => n9, ZN => n13);
   U14 : AOI222_X1 port map( A1 => B(9), A2 => n7, B1 => F(9), B2 => n5, C1 => 
                           C(9), C2 => n3, ZN => n12);
   U15 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => Y(8));
   U16 : AOI222_X1 port map( A1 => E(8), A2 => n11, B1 => A(8), B2 => n1, C1 =>
                           D(8), C2 => n9, ZN => n16);
   U17 : AOI222_X1 port map( A1 => B(8), A2 => n7, B1 => F(8), B2 => n5, C1 => 
                           C(8), C2 => n3, ZN => n15);
   U18 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => Y(7));
   U19 : AOI222_X1 port map( A1 => E(7), A2 => n11, B1 => A(7), B2 => n1, C1 =>
                           D(7), C2 => n9, ZN => n18);
   U20 : AOI222_X1 port map( A1 => B(7), A2 => n7, B1 => F(7), B2 => n5, C1 => 
                           C(7), C2 => n3, ZN => n17);
   U21 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => Y(6));
   U22 : AOI222_X1 port map( A1 => E(6), A2 => n11, B1 => A(6), B2 => n1, C1 =>
                           D(6), C2 => n9, ZN => n20);
   U23 : AOI222_X1 port map( A1 => B(6), A2 => n7, B1 => F(6), B2 => n5, C1 => 
                           C(6), C2 => n3, ZN => n19);
   U24 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => Y(5));
   U25 : AOI222_X1 port map( A1 => E(5), A2 => n11, B1 => A(5), B2 => n1, C1 =>
                           D(5), C2 => n9, ZN => n22);
   U26 : AOI222_X1 port map( A1 => B(5), A2 => n7, B1 => F(5), B2 => n5, C1 => 
                           C(5), C2 => n3, ZN => n21);
   U27 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => Y(4));
   U28 : AOI222_X1 port map( A1 => E(4), A2 => n11, B1 => A(4), B2 => n1, C1 =>
                           D(4), C2 => n9, ZN => n24);
   U29 : AOI222_X1 port map( A1 => B(4), A2 => n7, B1 => F(4), B2 => n5, C1 => 
                           C(4), C2 => n3, ZN => n23);
   U30 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => Y(3));
   U31 : AOI222_X1 port map( A1 => E(3), A2 => n11, B1 => A(3), B2 => n1, C1 =>
                           D(3), C2 => n9, ZN => n26);
   U32 : AOI222_X1 port map( A1 => B(3), A2 => n7, B1 => F(3), B2 => n5, C1 => 
                           C(3), C2 => n3, ZN => n25);
   U33 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => Y(31));
   U34 : AOI222_X1 port map( A1 => E(31), A2 => n11, B1 => A(31), B2 => n1, C1 
                           => D(31), C2 => n9, ZN => n28);
   U35 : AOI222_X1 port map( A1 => B(31), A2 => n7, B1 => F(31), B2 => n5, C1 
                           => C(31), C2 => n3, ZN => n27);
   U36 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => Y(30));
   U37 : AOI222_X1 port map( A1 => E(30), A2 => n11, B1 => A(30), B2 => n1, C1 
                           => D(30), C2 => n9, ZN => n30);
   U38 : AOI222_X1 port map( A1 => B(30), A2 => n7, B1 => F(30), B2 => n5, C1 
                           => C(30), C2 => n3, ZN => n29);
   U39 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => Y(2));
   U40 : AOI222_X1 port map( A1 => E(2), A2 => n11, B1 => A(2), B2 => n1, C1 =>
                           D(2), C2 => n9, ZN => n32);
   U41 : AOI222_X1 port map( A1 => B(2), A2 => n7, B1 => F(2), B2 => n5, C1 => 
                           C(2), C2 => n3, ZN => n31);
   U42 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => Y(29));
   U43 : AOI222_X1 port map( A1 => E(29), A2 => n11, B1 => A(29), B2 => n1, C1 
                           => D(29), C2 => n9, ZN => n34);
   U44 : AOI222_X1 port map( A1 => B(29), A2 => n7, B1 => F(29), B2 => n5, C1 
                           => C(29), C2 => n3, ZN => n33);
   U45 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => Y(28));
   U46 : AOI222_X1 port map( A1 => E(28), A2 => n11, B1 => A(28), B2 => n1, C1 
                           => D(28), C2 => n9, ZN => n36);
   U47 : AOI222_X1 port map( A1 => B(28), A2 => n7, B1 => F(28), B2 => n5, C1 
                           => C(28), C2 => n3, ZN => n35);
   U48 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => Y(27));
   U49 : AOI222_X1 port map( A1 => E(27), A2 => n11, B1 => A(27), B2 => n1, C1 
                           => D(27), C2 => n9, ZN => n38);
   U50 : AOI222_X1 port map( A1 => B(27), A2 => n7, B1 => F(27), B2 => n5, C1 
                           => C(27), C2 => n3, ZN => n37);
   U51 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => Y(26));
   U52 : AOI222_X1 port map( A1 => E(26), A2 => n11, B1 => A(26), B2 => n1, C1 
                           => D(26), C2 => n9, ZN => n40);
   U53 : AOI222_X1 port map( A1 => B(26), A2 => n7, B1 => F(26), B2 => n5, C1 
                           => C(26), C2 => n3, ZN => n39);
   U54 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => Y(25));
   U55 : AOI222_X1 port map( A1 => E(25), A2 => n11, B1 => A(25), B2 => n1, C1 
                           => D(25), C2 => n9, ZN => n42);
   U56 : AOI222_X1 port map( A1 => B(25), A2 => n7, B1 => F(25), B2 => n5, C1 
                           => C(25), C2 => n3, ZN => n41);
   U57 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => Y(24));
   U58 : AOI222_X1 port map( A1 => E(24), A2 => n11, B1 => A(24), B2 => n1, C1 
                           => D(24), C2 => n9, ZN => n44);
   U59 : AOI222_X1 port map( A1 => B(24), A2 => n7, B1 => F(24), B2 => n5, C1 
                           => C(24), C2 => n3, ZN => n43);
   U60 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => Y(23));
   U61 : AOI222_X1 port map( A1 => E(23), A2 => n11, B1 => A(23), B2 => n1, C1 
                           => D(23), C2 => n9, ZN => n46);
   U62 : AOI222_X1 port map( A1 => B(23), A2 => n7, B1 => F(23), B2 => n5, C1 
                           => C(23), C2 => n3, ZN => n45);
   U63 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => Y(22));
   U64 : AOI222_X1 port map( A1 => E(22), A2 => n11, B1 => A(22), B2 => n1, C1 
                           => D(22), C2 => n9, ZN => n48);
   U65 : AOI222_X1 port map( A1 => B(22), A2 => n7, B1 => F(22), B2 => n5, C1 
                           => C(22), C2 => n3, ZN => n47);
   U66 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => Y(21));
   U67 : AOI222_X1 port map( A1 => E(21), A2 => n11, B1 => A(21), B2 => n1, C1 
                           => D(21), C2 => n9, ZN => n50);
   U68 : AOI222_X1 port map( A1 => B(21), A2 => n7, B1 => F(21), B2 => n5, C1 
                           => C(21), C2 => n3, ZN => n49);
   U69 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => Y(20));
   U70 : AOI222_X1 port map( A1 => E(20), A2 => n11, B1 => A(20), B2 => n1, C1 
                           => D(20), C2 => n9, ZN => n52);
   U71 : AOI222_X1 port map( A1 => B(20), A2 => n7, B1 => F(20), B2 => n5, C1 
                           => C(20), C2 => n3, ZN => n51);
   U72 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => Y(1));
   U73 : AOI222_X1 port map( A1 => E(1), A2 => n11, B1 => A(1), B2 => n1, C1 =>
                           D(1), C2 => n9, ZN => n54);
   U74 : AOI222_X1 port map( A1 => B(1), A2 => n7, B1 => F(1), B2 => n5, C1 => 
                           C(1), C2 => n3, ZN => n53);
   U75 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => Y(19));
   U76 : AOI222_X1 port map( A1 => E(19), A2 => n11, B1 => A(19), B2 => n1, C1 
                           => D(19), C2 => n9, ZN => n56);
   U77 : AOI222_X1 port map( A1 => B(19), A2 => n7, B1 => F(19), B2 => n5, C1 
                           => C(19), C2 => n3, ZN => n55);
   U78 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => Y(18));
   U79 : AOI222_X1 port map( A1 => E(18), A2 => n11, B1 => A(18), B2 => n1, C1 
                           => D(18), C2 => n9, ZN => n58);
   U80 : AOI222_X1 port map( A1 => B(18), A2 => n7, B1 => F(18), B2 => n5, C1 
                           => C(18), C2 => n3, ZN => n57);
   U81 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => Y(17));
   U82 : AOI222_X1 port map( A1 => E(17), A2 => n11, B1 => A(17), B2 => n1, C1 
                           => D(17), C2 => n9, ZN => n60);
   U83 : AOI222_X1 port map( A1 => B(17), A2 => n7, B1 => F(17), B2 => n5, C1 
                           => C(17), C2 => n3, ZN => n59);
   U84 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => Y(16));
   U85 : AOI222_X1 port map( A1 => E(16), A2 => n11, B1 => A(16), B2 => n1, C1 
                           => D(16), C2 => n9, ZN => n62);
   U86 : AOI222_X1 port map( A1 => B(16), A2 => n7, B1 => F(16), B2 => n5, C1 
                           => C(16), C2 => n3, ZN => n61);
   U87 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => Y(15));
   U88 : AOI222_X1 port map( A1 => E(15), A2 => n11, B1 => A(15), B2 => n1, C1 
                           => D(15), C2 => n9, ZN => n64);
   U89 : AOI222_X1 port map( A1 => B(15), A2 => n7, B1 => F(15), B2 => n5, C1 
                           => C(15), C2 => n3, ZN => n63);
   U90 : NAND2_X1 port map( A1 => n65, A2 => n66, ZN => Y(14));
   U91 : AOI222_X1 port map( A1 => E(14), A2 => n11, B1 => A(14), B2 => n1, C1 
                           => D(14), C2 => n9, ZN => n66);
   U92 : AOI222_X1 port map( A1 => B(14), A2 => n7, B1 => F(14), B2 => n5, C1 
                           => C(14), C2 => n3, ZN => n65);
   U93 : NAND2_X1 port map( A1 => n67, A2 => n68, ZN => Y(13));
   U94 : AOI222_X1 port map( A1 => E(13), A2 => n11, B1 => A(13), B2 => n1, C1 
                           => D(13), C2 => n9, ZN => n68);
   U95 : AOI222_X1 port map( A1 => B(13), A2 => n7, B1 => F(13), B2 => n5, C1 
                           => C(13), C2 => n3, ZN => n67);
   U96 : NAND2_X1 port map( A1 => n69, A2 => n70, ZN => Y(12));
   U97 : AOI222_X1 port map( A1 => E(12), A2 => n11, B1 => A(12), B2 => n1, C1 
                           => D(12), C2 => n9, ZN => n70);
   U98 : AOI222_X1 port map( A1 => B(12), A2 => n7, B1 => F(12), B2 => n5, C1 
                           => C(12), C2 => n3, ZN => n69);
   U99 : NAND2_X1 port map( A1 => n71, A2 => n72, ZN => Y(11));
   U100 : AOI222_X1 port map( A1 => E(11), A2 => n11, B1 => A(11), B2 => n1, C1
                           => D(11), C2 => n9, ZN => n72);
   U101 : AOI222_X1 port map( A1 => B(11), A2 => n7, B1 => F(11), B2 => n5, C1 
                           => C(11), C2 => n3, ZN => n71);
   U102 : NAND2_X1 port map( A1 => n73, A2 => n74, ZN => Y(10));
   U103 : AOI222_X1 port map( A1 => E(10), A2 => n11, B1 => A(10), B2 => n1, C1
                           => D(10), C2 => n9, ZN => n74);
   U104 : AOI222_X1 port map( A1 => B(10), A2 => n7, B1 => F(10), B2 => n5, C1 
                           => C(10), C2 => n3, ZN => n73);
   U105 : NAND2_X1 port map( A1 => n75, A2 => n76, ZN => Y(0));
   U106 : AOI222_X1 port map( A1 => E(0), A2 => n11, B1 => A(0), B2 => n1, C1 
                           => D(0), C2 => n9, ZN => n76);
   U107 : NOR4_X1 port map( A1 => n9, A2 => n11, A3 => n77, A4 => n5, ZN => n14
                           );
   U108 : OR2_X1 port map( A1 => n7, A2 => n3, ZN => n77);
   U109 : AOI222_X1 port map( A1 => B(0), A2 => n7, B1 => F(0), B2 => n5, C1 =>
                           C(0), C2 => n3, ZN => n75);
   U110 : INV_X1 port map( A => S(1), ZN => n79);
   U111 : INV_X1 port map( A => S(2), ZN => n80);
   U112 : INV_X1 port map( A => S(0), ZN => n78);

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity MUX_2to1_n32 is

   port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : out 
         std_logic_vector (31 downto 0));

end MUX_2to1_n32;

architecture SYN_BEH of MUX_2to1_n32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(7), B => B(7), S => S, Z => Y(7));
   U2 : MUX2_X1 port map( A => A(6), B => B(6), S => S, Z => Y(6));
   U3 : MUX2_X1 port map( A => A(5), B => B(5), S => S, Z => Y(5));
   U4 : MUX2_X1 port map( A => A(4), B => B(4), S => S, Z => Y(4));
   U5 : MUX2_X1 port map( A => A(3), B => B(3), S => S, Z => Y(3));
   U6 : MUX2_X1 port map( A => A(2), B => B(2), S => S, Z => Y(2));
   U7 : MUX2_X1 port map( A => A(31), B => B(31), S => S, Z => Y(31));
   U8 : MUX2_X1 port map( A => A(30), B => B(30), S => S, Z => Y(30));
   U9 : MUX2_X1 port map( A => A(29), B => B(29), S => S, Z => Y(29));
   U10 : MUX2_X1 port map( A => A(28), B => B(28), S => S, Z => Y(28));
   U11 : MUX2_X1 port map( A => A(1), B => B(1), S => S, Z => Y(1));
   U12 : MUX2_X1 port map( A => A(27), B => B(27), S => S, Z => Y(27));
   U13 : MUX2_X1 port map( A => A(26), B => B(26), S => S, Z => Y(26));
   U14 : MUX2_X1 port map( A => A(25), B => B(25), S => S, Z => Y(25));
   U15 : MUX2_X1 port map( A => A(24), B => B(24), S => S, Z => Y(24));
   U16 : MUX2_X1 port map( A => A(23), B => B(23), S => S, Z => Y(23));
   U17 : MUX2_X1 port map( A => A(22), B => B(22), S => S, Z => Y(22));
   U18 : MUX2_X1 port map( A => A(21), B => B(21), S => S, Z => Y(21));
   U19 : MUX2_X1 port map( A => A(20), B => B(20), S => S, Z => Y(20));
   U20 : MUX2_X1 port map( A => A(19), B => B(19), S => S, Z => Y(19));
   U21 : MUX2_X1 port map( A => A(18), B => B(18), S => S, Z => Y(18));
   U22 : MUX2_X1 port map( A => A(0), B => B(0), S => S, Z => Y(0));
   U23 : MUX2_X1 port map( A => A(17), B => B(17), S => S, Z => Y(17));
   U24 : MUX2_X1 port map( A => A(16), B => B(16), S => S, Z => Y(16));
   U25 : MUX2_X1 port map( A => A(15), B => B(15), S => S, Z => Y(15));
   U26 : MUX2_X1 port map( A => A(14), B => B(14), S => S, Z => Y(14));
   U27 : MUX2_X1 port map( A => A(13), B => B(13), S => S, Z => Y(13));
   U28 : MUX2_X1 port map( A => A(12), B => B(12), S => S, Z => Y(12));
   U29 : MUX2_X1 port map( A => A(11), B => B(11), S => S, Z => Y(11));
   U30 : MUX2_X1 port map( A => A(10), B => B(10), S => S, Z => Y(10));
   U31 : MUX2_X1 port map( A => A(9), B => B(9), S => S, Z => Y(9));
   U32 : MUX2_X1 port map( A => A(8), B => B(8), S => S, Z => Y(8));

end SYN_BEH;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity compare_N32 is

   port( num1, num2 : in std_logic_vector (31 downto 0);  less, equal, greater 
         : out std_logic);

end compare_N32;

architecture SYN_Behavioral of compare_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   signal greater_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
      n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28
      , n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, 
      n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57
      , n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, 
      n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86
      , n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, 
      n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111 : 
      std_logic;

begin
   greater <= greater_port;
   
   U2 : AOI21_X1 port map( B1 => n1, B2 => n2, A => greater_port, ZN => less);
   U3 : INV_X1 port map( A => n3, ZN => n1);
   U4 : NOR3_X1 port map( A1 => n3, A2 => greater_port, A3 => n4, ZN => equal);
   U5 : INV_X1 port map( A => n2, ZN => n4);
   U6 : OAI22_X1 port map( A1 => n5, A2 => n6, B1 => num2(31), B2 => n7, ZN => 
                           greater_port);
   U7 : NAND2_X1 port map( A1 => n2, A2 => n8, ZN => n6);
   U8 : NAND2_X1 port map( A1 => num2(31), A2 => n7, ZN => n2);
   U9 : INV_X1 port map( A => num1(31), ZN => n7);
   U10 : AOI22_X1 port map( A1 => num1(30), A2 => n9, B1 => n10, B2 => n11, ZN 
                           => n5);
   U11 : OAI221_X1 port map( B1 => num2(29), B2 => n12, C1 => num2(28), C2 => 
                           n13, A => n14, ZN => n11);
   U12 : NAND3_X1 port map( A1 => n15, A2 => n16, A3 => n17, ZN => n14);
   U13 : OAI221_X1 port map( B1 => num2(27), B2 => n18, C1 => num2(26), C2 => 
                           n19, A => n20, ZN => n16);
   U14 : NAND3_X1 port map( A1 => n21, A2 => n22, A3 => n23, ZN => n20);
   U15 : OAI221_X1 port map( B1 => num2(25), B2 => n24, C1 => num2(24), C2 => 
                           n25, A => n26, ZN => n22);
   U16 : NAND3_X1 port map( A1 => n27, A2 => n28, A3 => n29, ZN => n26);
   U17 : OAI221_X1 port map( B1 => num2(23), B2 => n30, C1 => num2(22), C2 => 
                           n31, A => n32, ZN => n28);
   U18 : NAND3_X1 port map( A1 => n33, A2 => n34, A3 => n35, ZN => n32);
   U19 : OAI221_X1 port map( B1 => num2(21), B2 => n36, C1 => num2(20), C2 => 
                           n37, A => n38, ZN => n34);
   U20 : NAND3_X1 port map( A1 => n39, A2 => n40, A3 => n41, ZN => n38);
   U21 : OAI221_X1 port map( B1 => num2(19), B2 => n42, C1 => num2(18), C2 => 
                           n43, A => n44, ZN => n40);
   U22 : NAND3_X1 port map( A1 => n45, A2 => n46, A3 => n47, ZN => n44);
   U23 : OAI221_X1 port map( B1 => num2(17), B2 => n48, C1 => num2(16), C2 => 
                           n49, A => n50, ZN => n46);
   U24 : NAND3_X1 port map( A1 => n51, A2 => n52, A3 => n53, ZN => n50);
   U25 : OAI221_X1 port map( B1 => num2(15), B2 => n54, C1 => num2(14), C2 => 
                           n55, A => n56, ZN => n52);
   U26 : NAND3_X1 port map( A1 => n57, A2 => n58, A3 => n59, ZN => n56);
   U27 : OAI221_X1 port map( B1 => num2(13), B2 => n60, C1 => num2(12), C2 => 
                           n61, A => n62, ZN => n58);
   U28 : NAND3_X1 port map( A1 => n63, A2 => n64, A3 => n65, ZN => n62);
   U29 : OAI221_X1 port map( B1 => num2(11), B2 => n66, C1 => num2(10), C2 => 
                           n67, A => n68, ZN => n64);
   U30 : NAND3_X1 port map( A1 => n69, A2 => n70, A3 => n71, ZN => n68);
   U31 : OAI221_X1 port map( B1 => num2(9), B2 => n72, C1 => num2(8), C2 => n73
                           , A => n74, ZN => n70);
   U32 : NAND3_X1 port map( A1 => n75, A2 => n76, A3 => n77, ZN => n74);
   U33 : OAI221_X1 port map( B1 => num2(7), B2 => n78, C1 => num2(6), C2 => n79
                           , A => n80, ZN => n76);
   U34 : NAND3_X1 port map( A1 => n81, A2 => n82, A3 => n83, ZN => n80);
   U35 : OAI221_X1 port map( B1 => num2(5), B2 => n84, C1 => num2(4), C2 => n85
                           , A => n86, ZN => n82);
   U36 : NAND3_X1 port map( A1 => n87, A2 => n88, A3 => n89, ZN => n86);
   U37 : OAI221_X1 port map( B1 => num2(3), B2 => n90, C1 => num2(2), C2 => n91
                           , A => n92, ZN => n88);
   U38 : OAI211_X1 port map( C1 => num1(1), C2 => n93, A => n94, B => n95, ZN 
                           => n92);
   U39 : OAI21_X1 port map( B1 => num2(0), B2 => n96, A => num2(1), ZN => n95);
   U40 : NOR3_X1 port map( A1 => n96, A2 => num2(1), A3 => num2(0), ZN => n93);
   U41 : NAND3_X1 port map( A1 => n97, A2 => n98, A3 => n99, ZN => n3);
   U42 : NOR4_X1 port map( A1 => n100, A2 => n101, A3 => n102, A4 => n103, ZN 
                           => n99);
   U43 : NAND3_X1 port map( A1 => n17, A2 => n15, A3 => n10, ZN => n103);
   U44 : NAND2_X1 port map( A1 => num2(29), A2 => n12, ZN => n10);
   U45 : INV_X1 port map( A => num1(29), ZN => n12);
   U46 : NAND2_X1 port map( A1 => num2(28), A2 => n13, ZN => n15);
   U47 : INV_X1 port map( A => num1(28), ZN => n13);
   U48 : NAND2_X1 port map( A1 => num2(27), A2 => n18, ZN => n17);
   U49 : INV_X1 port map( A => num1(27), ZN => n18);
   U50 : NAND4_X1 port map( A1 => n23, A2 => n21, A3 => n29, A4 => n27, ZN => 
                           n102);
   U51 : NAND2_X1 port map( A1 => num2(24), A2 => n25, ZN => n27);
   U52 : INV_X1 port map( A => num1(24), ZN => n25);
   U53 : NAND2_X1 port map( A1 => num2(23), A2 => n30, ZN => n29);
   U54 : INV_X1 port map( A => num1(23), ZN => n30);
   U55 : NAND2_X1 port map( A1 => num2(26), A2 => n19, ZN => n21);
   U56 : INV_X1 port map( A => num1(26), ZN => n19);
   U57 : NAND2_X1 port map( A1 => num2(25), A2 => n24, ZN => n23);
   U58 : INV_X1 port map( A => num1(25), ZN => n24);
   U59 : NAND4_X1 port map( A1 => n35, A2 => n33, A3 => n41, A4 => n39, ZN => 
                           n101);
   U60 : NAND2_X1 port map( A1 => num2(20), A2 => n37, ZN => n39);
   U61 : INV_X1 port map( A => num1(20), ZN => n37);
   U62 : NAND2_X1 port map( A1 => num2(19), A2 => n42, ZN => n41);
   U63 : INV_X1 port map( A => num1(19), ZN => n42);
   U64 : NAND2_X1 port map( A1 => num2(22), A2 => n31, ZN => n33);
   U65 : INV_X1 port map( A => num1(22), ZN => n31);
   U66 : NAND2_X1 port map( A1 => num2(21), A2 => n36, ZN => n35);
   U67 : INV_X1 port map( A => num1(21), ZN => n36);
   U68 : NAND4_X1 port map( A1 => n47, A2 => n45, A3 => n53, A4 => n51, ZN => 
                           n100);
   U69 : NAND2_X1 port map( A1 => num2(16), A2 => n49, ZN => n51);
   U70 : INV_X1 port map( A => num1(16), ZN => n49);
   U71 : NAND2_X1 port map( A1 => num2(15), A2 => n54, ZN => n53);
   U72 : INV_X1 port map( A => num1(15), ZN => n54);
   U73 : NAND2_X1 port map( A1 => num2(18), A2 => n43, ZN => n45);
   U74 : INV_X1 port map( A => num1(18), ZN => n43);
   U75 : NAND2_X1 port map( A1 => num2(17), A2 => n48, ZN => n47);
   U76 : INV_X1 port map( A => num1(17), ZN => n48);
   U77 : NOR4_X1 port map( A1 => n104, A2 => n105, A3 => n106, A4 => n107, ZN 
                           => n98);
   U78 : INV_X1 port map( A => n87, ZN => n107);
   U79 : NAND2_X1 port map( A1 => num2(4), A2 => n85, ZN => n87);
   U80 : INV_X1 port map( A => num1(4), ZN => n85);
   U81 : INV_X1 port map( A => n94, ZN => n106);
   U82 : NAND2_X1 port map( A1 => num2(2), A2 => n91, ZN => n94);
   U83 : INV_X1 port map( A => num1(2), ZN => n91);
   U84 : OAI21_X1 port map( B1 => n108, B2 => n109, A => n8, ZN => n105);
   U85 : OR2_X1 port map( A1 => n9, A2 => num1(30), ZN => n8);
   U86 : INV_X1 port map( A => num2(30), ZN => n9);
   U87 : AOI21_X1 port map( B1 => num2(0), B2 => n96, A => n110, ZN => n109);
   U88 : INV_X1 port map( A => num1(1), ZN => n110);
   U89 : AOI21_X1 port map( B1 => num2(0), B2 => n96, A => num2(1), ZN => n108)
                           ;
   U90 : INV_X1 port map( A => num1(0), ZN => n96);
   U91 : NAND4_X1 port map( A1 => n75, A2 => n83, A3 => n81, A4 => n89, ZN => 
                           n104);
   U92 : NAND2_X1 port map( A1 => num2(3), A2 => n90, ZN => n89);
   U93 : INV_X1 port map( A => num1(3), ZN => n90);
   U94 : NAND2_X1 port map( A1 => num2(6), A2 => n79, ZN => n81);
   U95 : INV_X1 port map( A => num1(6), ZN => n79);
   U96 : NAND2_X1 port map( A1 => num2(5), A2 => n84, ZN => n83);
   U97 : INV_X1 port map( A => num1(5), ZN => n84);
   U98 : NAND2_X1 port map( A1 => num2(8), A2 => n73, ZN => n75);
   U99 : INV_X1 port map( A => num1(8), ZN => n73);
   U100 : AND4_X1 port map( A1 => n111, A2 => n59, A3 => n65, A4 => n57, ZN => 
                           n97);
   U101 : NAND2_X1 port map( A1 => num2(14), A2 => n55, ZN => n57);
   U102 : INV_X1 port map( A => num1(14), ZN => n55);
   U103 : NAND2_X1 port map( A1 => num2(11), A2 => n66, ZN => n65);
   U104 : INV_X1 port map( A => num1(11), ZN => n66);
   U105 : NAND2_X1 port map( A1 => num2(13), A2 => n60, ZN => n59);
   U106 : INV_X1 port map( A => num1(13), ZN => n60);
   U107 : AND4_X1 port map( A1 => n63, A2 => n71, A3 => n69, A4 => n77, ZN => 
                           n111);
   U108 : NAND2_X1 port map( A1 => num2(7), A2 => n78, ZN => n77);
   U109 : INV_X1 port map( A => num1(7), ZN => n78);
   U110 : NAND2_X1 port map( A1 => num2(9), A2 => n72, ZN => n69);
   U111 : INV_X1 port map( A => num1(9), ZN => n72);
   U112 : NAND2_X1 port map( A1 => num2(10), A2 => n67, ZN => n71);
   U113 : INV_X1 port map( A => num1(10), ZN => n67);
   U114 : NAND2_X1 port map( A1 => num2(12), A2 => n61, ZN => n63);
   U115 : INV_X1 port map( A => num1(12), ZN => n61);

end SYN_Behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity p4_adder_N32_N_carry4 is

   port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  SUM : 
         out std_logic_vector (31 downto 0));

end p4_adder_N32_N_carry4;

architecture SYN_beh of p4_adder_N32_N_carry4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component sum_generator_N32_N_carry4
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic_vector
            (8 downto 0);  Sum : out std_logic_vector (31 downto 0));
   end component;
   
   component sparse_tree_carry_gen_N5
      port( A, B : in std_logic_vector (31 downto 0);  C0 : in std_logic;  Cout
            : out std_logic_vector (7 downto 0));
   end component;
   
   signal notb_31_port, notb_30_port, notb_29_port, notb_28_port, notb_27_port,
      notb_26_port, notb_25_port, notb_24_port, notb_23_port, notb_22_port, 
      notb_21_port, notb_20_port, notb_19_port, notb_18_port, notb_17_port, 
      notb_16_port, notb_15_port, notb_14_port, notb_13_port, notb_12_port, 
      notb_11_port, notb_10_port, notb_9_port, notb_8_port, notb_7_port, 
      notb_6_port, notb_5_port, notb_4_port, notb_3_port, notb_2_port, 
      notb_1_port, notb_0_port, carry_7_port, carry_6_port, carry_5_port, 
      carry_4_port, carry_3_port, carry_2_port, carry_1_port, carry_0_port : 
      std_logic;

begin
   
   sparsetree : sparse_tree_carry_gen_N5 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), B(31) => notb_31_port, B(30) 
                           => notb_30_port, B(29) => notb_29_port, B(28) => 
                           notb_28_port, B(27) => notb_27_port, B(26) => 
                           notb_26_port, B(25) => notb_25_port, B(24) => 
                           notb_24_port, B(23) => notb_23_port, B(22) => 
                           notb_22_port, B(21) => notb_21_port, B(20) => 
                           notb_20_port, B(19) => notb_19_port, B(18) => 
                           notb_18_port, B(17) => notb_17_port, B(16) => 
                           notb_16_port, B(15) => notb_15_port, B(14) => 
                           notb_14_port, B(13) => notb_13_port, B(12) => 
                           notb_12_port, B(11) => notb_11_port, B(10) => 
                           notb_10_port, B(9) => notb_9_port, B(8) => 
                           notb_8_port, B(7) => notb_7_port, B(6) => 
                           notb_6_port, B(5) => notb_5_port, B(4) => 
                           notb_4_port, B(3) => notb_3_port, B(2) => 
                           notb_2_port, B(1) => notb_1_port, B(0) => 
                           notb_0_port, C0 => Cin, Cout(7) => carry_7_port, 
                           Cout(6) => carry_6_port, Cout(5) => carry_5_port, 
                           Cout(4) => carry_4_port, Cout(3) => carry_3_port, 
                           Cout(2) => carry_2_port, Cout(1) => carry_1_port, 
                           Cout(0) => carry_0_port);
   sumgen : sum_generator_N32_N_carry4 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), B(31) => notb_31_port, B(30) => 
                           notb_30_port, B(29) => notb_29_port, B(28) => 
                           notb_28_port, B(27) => notb_27_port, B(26) => 
                           notb_26_port, B(25) => notb_25_port, B(24) => 
                           notb_24_port, B(23) => notb_23_port, B(22) => 
                           notb_22_port, B(21) => notb_21_port, B(20) => 
                           notb_20_port, B(19) => notb_19_port, B(18) => 
                           notb_18_port, B(17) => notb_17_port, B(16) => 
                           notb_16_port, B(15) => notb_15_port, B(14) => 
                           notb_14_port, B(13) => notb_13_port, B(12) => 
                           notb_12_port, B(11) => notb_11_port, B(10) => 
                           notb_10_port, B(9) => notb_9_port, B(8) => 
                           notb_8_port, B(7) => notb_7_port, B(6) => 
                           notb_6_port, B(5) => notb_5_port, B(4) => 
                           notb_4_port, B(3) => notb_3_port, B(2) => 
                           notb_2_port, B(1) => notb_1_port, B(0) => 
                           notb_0_port, Ci(8) => carry_7_port, Ci(7) => 
                           carry_6_port, Ci(6) => carry_5_port, Ci(5) => 
                           carry_4_port, Ci(4) => carry_3_port, Ci(3) => 
                           carry_2_port, Ci(2) => carry_1_port, Ci(1) => 
                           carry_0_port, Ci(0) => Cin, Sum(31) => SUM(31), 
                           Sum(30) => SUM(30), Sum(29) => SUM(29), Sum(28) => 
                           SUM(28), Sum(27) => SUM(27), Sum(26) => SUM(26), 
                           Sum(25) => SUM(25), Sum(24) => SUM(24), Sum(23) => 
                           SUM(23), Sum(22) => SUM(22), Sum(21) => SUM(21), 
                           Sum(20) => SUM(20), Sum(19) => SUM(19), Sum(18) => 
                           SUM(18), Sum(17) => SUM(17), Sum(16) => SUM(16), 
                           Sum(15) => SUM(15), Sum(14) => SUM(14), Sum(13) => 
                           SUM(13), Sum(12) => SUM(12), Sum(11) => SUM(11), 
                           Sum(10) => SUM(10), Sum(9) => SUM(9), Sum(8) => 
                           SUM(8), Sum(7) => SUM(7), Sum(6) => SUM(6), Sum(5) 
                           => SUM(5), Sum(4) => SUM(4), Sum(3) => SUM(3), 
                           Sum(2) => SUM(2), Sum(1) => SUM(1), Sum(0) => SUM(0)
                           );
   U1 : XOR2_X1 port map( A => Cin, B => B(9), Z => notb_9_port);
   U2 : XOR2_X1 port map( A => Cin, B => B(8), Z => notb_8_port);
   U3 : XOR2_X1 port map( A => Cin, B => B(7), Z => notb_7_port);
   U4 : XOR2_X1 port map( A => Cin, B => B(6), Z => notb_6_port);
   U5 : XOR2_X1 port map( A => Cin, B => B(5), Z => notb_5_port);
   U6 : XOR2_X1 port map( A => Cin, B => B(4), Z => notb_4_port);
   U7 : XOR2_X1 port map( A => Cin, B => B(3), Z => notb_3_port);
   U8 : XOR2_X1 port map( A => Cin, B => B(31), Z => notb_31_port);
   U9 : XOR2_X1 port map( A => Cin, B => B(30), Z => notb_30_port);
   U10 : XOR2_X1 port map( A => Cin, B => B(2), Z => notb_2_port);
   U11 : XOR2_X1 port map( A => Cin, B => B(29), Z => notb_29_port);
   U12 : XOR2_X1 port map( A => Cin, B => B(28), Z => notb_28_port);
   U13 : XOR2_X1 port map( A => Cin, B => B(27), Z => notb_27_port);
   U14 : XOR2_X1 port map( A => Cin, B => B(26), Z => notb_26_port);
   U15 : XOR2_X1 port map( A => Cin, B => B(25), Z => notb_25_port);
   U16 : XOR2_X1 port map( A => Cin, B => B(24), Z => notb_24_port);
   U17 : XOR2_X1 port map( A => Cin, B => B(23), Z => notb_23_port);
   U18 : XOR2_X1 port map( A => Cin, B => B(22), Z => notb_22_port);
   U19 : XOR2_X1 port map( A => Cin, B => B(21), Z => notb_21_port);
   U20 : XOR2_X1 port map( A => Cin, B => B(20), Z => notb_20_port);
   U21 : XOR2_X1 port map( A => Cin, B => B(1), Z => notb_1_port);
   U22 : XOR2_X1 port map( A => Cin, B => B(19), Z => notb_19_port);
   U23 : XOR2_X1 port map( A => Cin, B => B(18), Z => notb_18_port);
   U24 : XOR2_X1 port map( A => Cin, B => B(17), Z => notb_17_port);
   U25 : XOR2_X1 port map( A => Cin, B => B(16), Z => notb_16_port);
   U26 : XOR2_X1 port map( A => Cin, B => B(15), Z => notb_15_port);
   U27 : XOR2_X1 port map( A => Cin, B => B(14), Z => notb_14_port);
   U28 : XOR2_X1 port map( A => Cin, B => B(13), Z => notb_13_port);
   U29 : XOR2_X1 port map( A => Cin, B => B(12), Z => notb_12_port);
   U30 : XOR2_X1 port map( A => Cin, B => B(11), Z => notb_11_port);
   U31 : XOR2_X1 port map( A => Cin, B => B(10), Z => notb_10_port);
   U32 : XOR2_X1 port map( A => Cin, B => B(0), Z => notb_0_port);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity operatore_logic_REG_SIZE32 is

   port( A, B : in std_logic_vector (31 downto 0);  OUT_LOGIC_AND, OUT_LOGIC_OR
         , OUT_LOGIC_XOR : out std_logic_vector (31 downto 0));

end operatore_logic_REG_SIZE32;

architecture SYN_behaviour of operatore_logic_REG_SIZE32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   signal n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16
      , n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, 
      n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45
      , n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, 
      n60, n61, n62, n63, n64 : std_logic;

begin
   
   U1 : INV_X1 port map( A => B(4), ZN => n1);
   U2 : XOR2_X1 port map( A => B(9), B => A(9), Z => OUT_LOGIC_XOR(9));
   U3 : XOR2_X1 port map( A => B(8), B => A(8), Z => OUT_LOGIC_XOR(8));
   U4 : XOR2_X1 port map( A => B(7), B => A(7), Z => OUT_LOGIC_XOR(7));
   U5 : XOR2_X1 port map( A => B(6), B => A(6), Z => OUT_LOGIC_XOR(6));
   U6 : XOR2_X1 port map( A => B(5), B => A(5), Z => OUT_LOGIC_XOR(5));
   U7 : XOR2_X1 port map( A => B(4), B => A(4), Z => OUT_LOGIC_XOR(4));
   U8 : XOR2_X1 port map( A => B(3), B => A(3), Z => OUT_LOGIC_XOR(3));
   U9 : XOR2_X1 port map( A => B(31), B => A(31), Z => OUT_LOGIC_XOR(31));
   U10 : XOR2_X1 port map( A => B(30), B => A(30), Z => OUT_LOGIC_XOR(30));
   U11 : XOR2_X1 port map( A => B(2), B => A(2), Z => OUT_LOGIC_XOR(2));
   U12 : XOR2_X1 port map( A => B(29), B => A(29), Z => OUT_LOGIC_XOR(29));
   U13 : XOR2_X1 port map( A => B(28), B => A(28), Z => OUT_LOGIC_XOR(28));
   U14 : XOR2_X1 port map( A => B(27), B => A(27), Z => OUT_LOGIC_XOR(27));
   U15 : XOR2_X1 port map( A => B(26), B => A(26), Z => OUT_LOGIC_XOR(26));
   U16 : XOR2_X1 port map( A => B(25), B => A(25), Z => OUT_LOGIC_XOR(25));
   U17 : XOR2_X1 port map( A => B(24), B => A(24), Z => OUT_LOGIC_XOR(24));
   U18 : XOR2_X1 port map( A => B(23), B => A(23), Z => OUT_LOGIC_XOR(23));
   U19 : XOR2_X1 port map( A => B(22), B => A(22), Z => OUT_LOGIC_XOR(22));
   U20 : XOR2_X1 port map( A => B(21), B => A(21), Z => OUT_LOGIC_XOR(21));
   U21 : XOR2_X1 port map( A => B(20), B => A(20), Z => OUT_LOGIC_XOR(20));
   U22 : XOR2_X1 port map( A => B(1), B => A(1), Z => OUT_LOGIC_XOR(1));
   U23 : XOR2_X1 port map( A => B(19), B => A(19), Z => OUT_LOGIC_XOR(19));
   U24 : XOR2_X1 port map( A => B(18), B => A(18), Z => OUT_LOGIC_XOR(18));
   U25 : XOR2_X1 port map( A => B(17), B => A(17), Z => OUT_LOGIC_XOR(17));
   U26 : XOR2_X1 port map( A => B(16), B => A(16), Z => OUT_LOGIC_XOR(16));
   U27 : XOR2_X1 port map( A => B(15), B => A(15), Z => OUT_LOGIC_XOR(15));
   U28 : XOR2_X1 port map( A => B(14), B => A(14), Z => OUT_LOGIC_XOR(14));
   U29 : XOR2_X1 port map( A => B(13), B => A(13), Z => OUT_LOGIC_XOR(13));
   U30 : XOR2_X1 port map( A => B(12), B => A(12), Z => OUT_LOGIC_XOR(12));
   U31 : XOR2_X1 port map( A => B(11), B => A(11), Z => OUT_LOGIC_XOR(11));
   U32 : XOR2_X1 port map( A => B(10), B => A(10), Z => OUT_LOGIC_XOR(10));
   U33 : XOR2_X1 port map( A => B(0), B => A(0), Z => OUT_LOGIC_XOR(0));
   U34 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => OUT_LOGIC_OR(9));
   U35 : NAND2_X1 port map( A1 => n4, A2 => n5, ZN => OUT_LOGIC_OR(8));
   U36 : NAND2_X1 port map( A1 => n6, A2 => n7, ZN => OUT_LOGIC_OR(7));
   U37 : NAND2_X1 port map( A1 => n8, A2 => n9, ZN => OUT_LOGIC_OR(6));
   U38 : NAND2_X1 port map( A1 => n10, A2 => n11, ZN => OUT_LOGIC_OR(5));
   U39 : NAND2_X1 port map( A1 => n1, A2 => n12, ZN => OUT_LOGIC_OR(4));
   U40 : NAND2_X1 port map( A1 => n13, A2 => n14, ZN => OUT_LOGIC_OR(3));
   U41 : NAND2_X1 port map( A1 => n15, A2 => n16, ZN => OUT_LOGIC_OR(31));
   U42 : NAND2_X1 port map( A1 => n17, A2 => n18, ZN => OUT_LOGIC_OR(30));
   U43 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => OUT_LOGIC_OR(2));
   U44 : NAND2_X1 port map( A1 => n21, A2 => n22, ZN => OUT_LOGIC_OR(29));
   U45 : NAND2_X1 port map( A1 => n23, A2 => n24, ZN => OUT_LOGIC_OR(28));
   U46 : NAND2_X1 port map( A1 => n25, A2 => n26, ZN => OUT_LOGIC_OR(27));
   U47 : NAND2_X1 port map( A1 => n27, A2 => n28, ZN => OUT_LOGIC_OR(26));
   U48 : NAND2_X1 port map( A1 => n29, A2 => n30, ZN => OUT_LOGIC_OR(25));
   U49 : NAND2_X1 port map( A1 => n31, A2 => n32, ZN => OUT_LOGIC_OR(24));
   U50 : NAND2_X1 port map( A1 => n33, A2 => n34, ZN => OUT_LOGIC_OR(23));
   U51 : NAND2_X1 port map( A1 => n35, A2 => n36, ZN => OUT_LOGIC_OR(22));
   U52 : NAND2_X1 port map( A1 => n37, A2 => n38, ZN => OUT_LOGIC_OR(21));
   U53 : NAND2_X1 port map( A1 => n39, A2 => n40, ZN => OUT_LOGIC_OR(20));
   U54 : NAND2_X1 port map( A1 => n41, A2 => n42, ZN => OUT_LOGIC_OR(1));
   U55 : NAND2_X1 port map( A1 => n43, A2 => n44, ZN => OUT_LOGIC_OR(19));
   U56 : NAND2_X1 port map( A1 => n45, A2 => n46, ZN => OUT_LOGIC_OR(18));
   U57 : NAND2_X1 port map( A1 => n47, A2 => n48, ZN => OUT_LOGIC_OR(17));
   U58 : NAND2_X1 port map( A1 => n49, A2 => n50, ZN => OUT_LOGIC_OR(16));
   U59 : NAND2_X1 port map( A1 => n51, A2 => n52, ZN => OUT_LOGIC_OR(15));
   U60 : NAND2_X1 port map( A1 => n53, A2 => n54, ZN => OUT_LOGIC_OR(14));
   U61 : NAND2_X1 port map( A1 => n55, A2 => n56, ZN => OUT_LOGIC_OR(13));
   U62 : NAND2_X1 port map( A1 => n57, A2 => n58, ZN => OUT_LOGIC_OR(12));
   U63 : NAND2_X1 port map( A1 => n59, A2 => n60, ZN => OUT_LOGIC_OR(11));
   U64 : NAND2_X1 port map( A1 => n61, A2 => n62, ZN => OUT_LOGIC_OR(10));
   U65 : NAND2_X1 port map( A1 => n63, A2 => n64, ZN => OUT_LOGIC_OR(0));
   U66 : NOR2_X1 port map( A1 => n2, A2 => n3, ZN => OUT_LOGIC_AND(9));
   U67 : INV_X1 port map( A => A(9), ZN => n3);
   U68 : INV_X1 port map( A => B(9), ZN => n2);
   U69 : NOR2_X1 port map( A1 => n4, A2 => n5, ZN => OUT_LOGIC_AND(8));
   U70 : INV_X1 port map( A => A(8), ZN => n5);
   U71 : INV_X1 port map( A => B(8), ZN => n4);
   U72 : NOR2_X1 port map( A1 => n6, A2 => n7, ZN => OUT_LOGIC_AND(7));
   U73 : INV_X1 port map( A => A(7), ZN => n7);
   U74 : INV_X1 port map( A => B(7), ZN => n6);
   U75 : NOR2_X1 port map( A1 => n8, A2 => n9, ZN => OUT_LOGIC_AND(6));
   U76 : INV_X1 port map( A => A(6), ZN => n9);
   U77 : INV_X1 port map( A => B(6), ZN => n8);
   U78 : NOR2_X1 port map( A1 => n10, A2 => n11, ZN => OUT_LOGIC_AND(5));
   U79 : INV_X1 port map( A => A(5), ZN => n11);
   U80 : INV_X1 port map( A => B(5), ZN => n10);
   U81 : NOR2_X1 port map( A1 => n1, A2 => n12, ZN => OUT_LOGIC_AND(4));
   U82 : INV_X1 port map( A => A(4), ZN => n12);
   U83 : NOR2_X1 port map( A1 => n13, A2 => n14, ZN => OUT_LOGIC_AND(3));
   U84 : INV_X1 port map( A => A(3), ZN => n14);
   U85 : INV_X1 port map( A => B(3), ZN => n13);
   U86 : NOR2_X1 port map( A1 => n15, A2 => n16, ZN => OUT_LOGIC_AND(31));
   U87 : INV_X1 port map( A => A(31), ZN => n16);
   U88 : INV_X1 port map( A => B(31), ZN => n15);
   U89 : NOR2_X1 port map( A1 => n17, A2 => n18, ZN => OUT_LOGIC_AND(30));
   U90 : INV_X1 port map( A => A(30), ZN => n18);
   U91 : INV_X1 port map( A => B(30), ZN => n17);
   U92 : NOR2_X1 port map( A1 => n19, A2 => n20, ZN => OUT_LOGIC_AND(2));
   U93 : INV_X1 port map( A => A(2), ZN => n20);
   U94 : INV_X1 port map( A => B(2), ZN => n19);
   U95 : NOR2_X1 port map( A1 => n21, A2 => n22, ZN => OUT_LOGIC_AND(29));
   U96 : INV_X1 port map( A => A(29), ZN => n22);
   U97 : INV_X1 port map( A => B(29), ZN => n21);
   U98 : NOR2_X1 port map( A1 => n23, A2 => n24, ZN => OUT_LOGIC_AND(28));
   U99 : INV_X1 port map( A => A(28), ZN => n24);
   U100 : INV_X1 port map( A => B(28), ZN => n23);
   U101 : NOR2_X1 port map( A1 => n25, A2 => n26, ZN => OUT_LOGIC_AND(27));
   U102 : INV_X1 port map( A => A(27), ZN => n26);
   U103 : INV_X1 port map( A => B(27), ZN => n25);
   U104 : NOR2_X1 port map( A1 => n27, A2 => n28, ZN => OUT_LOGIC_AND(26));
   U105 : INV_X1 port map( A => A(26), ZN => n28);
   U106 : INV_X1 port map( A => B(26), ZN => n27);
   U107 : NOR2_X1 port map( A1 => n29, A2 => n30, ZN => OUT_LOGIC_AND(25));
   U108 : INV_X1 port map( A => A(25), ZN => n30);
   U109 : INV_X1 port map( A => B(25), ZN => n29);
   U110 : NOR2_X1 port map( A1 => n31, A2 => n32, ZN => OUT_LOGIC_AND(24));
   U111 : INV_X1 port map( A => A(24), ZN => n32);
   U112 : INV_X1 port map( A => B(24), ZN => n31);
   U113 : NOR2_X1 port map( A1 => n33, A2 => n34, ZN => OUT_LOGIC_AND(23));
   U114 : INV_X1 port map( A => A(23), ZN => n34);
   U115 : INV_X1 port map( A => B(23), ZN => n33);
   U116 : NOR2_X1 port map( A1 => n35, A2 => n36, ZN => OUT_LOGIC_AND(22));
   U117 : INV_X1 port map( A => A(22), ZN => n36);
   U118 : INV_X1 port map( A => B(22), ZN => n35);
   U119 : NOR2_X1 port map( A1 => n37, A2 => n38, ZN => OUT_LOGIC_AND(21));
   U120 : INV_X1 port map( A => A(21), ZN => n38);
   U121 : INV_X1 port map( A => B(21), ZN => n37);
   U122 : NOR2_X1 port map( A1 => n39, A2 => n40, ZN => OUT_LOGIC_AND(20));
   U123 : INV_X1 port map( A => A(20), ZN => n40);
   U124 : INV_X1 port map( A => B(20), ZN => n39);
   U125 : NOR2_X1 port map( A1 => n41, A2 => n42, ZN => OUT_LOGIC_AND(1));
   U126 : INV_X1 port map( A => A(1), ZN => n42);
   U127 : INV_X1 port map( A => B(1), ZN => n41);
   U128 : NOR2_X1 port map( A1 => n43, A2 => n44, ZN => OUT_LOGIC_AND(19));
   U129 : INV_X1 port map( A => A(19), ZN => n44);
   U130 : INV_X1 port map( A => B(19), ZN => n43);
   U131 : NOR2_X1 port map( A1 => n45, A2 => n46, ZN => OUT_LOGIC_AND(18));
   U132 : INV_X1 port map( A => A(18), ZN => n46);
   U133 : INV_X1 port map( A => B(18), ZN => n45);
   U134 : NOR2_X1 port map( A1 => n47, A2 => n48, ZN => OUT_LOGIC_AND(17));
   U135 : INV_X1 port map( A => A(17), ZN => n48);
   U136 : INV_X1 port map( A => B(17), ZN => n47);
   U137 : NOR2_X1 port map( A1 => n49, A2 => n50, ZN => OUT_LOGIC_AND(16));
   U138 : INV_X1 port map( A => A(16), ZN => n50);
   U139 : INV_X1 port map( A => B(16), ZN => n49);
   U140 : NOR2_X1 port map( A1 => n51, A2 => n52, ZN => OUT_LOGIC_AND(15));
   U141 : INV_X1 port map( A => A(15), ZN => n52);
   U142 : INV_X1 port map( A => B(15), ZN => n51);
   U143 : NOR2_X1 port map( A1 => n53, A2 => n54, ZN => OUT_LOGIC_AND(14));
   U144 : INV_X1 port map( A => A(14), ZN => n54);
   U145 : INV_X1 port map( A => B(14), ZN => n53);
   U146 : NOR2_X1 port map( A1 => n55, A2 => n56, ZN => OUT_LOGIC_AND(13));
   U147 : INV_X1 port map( A => A(13), ZN => n56);
   U148 : INV_X1 port map( A => B(13), ZN => n55);
   U149 : NOR2_X1 port map( A1 => n57, A2 => n58, ZN => OUT_LOGIC_AND(12));
   U150 : INV_X1 port map( A => A(12), ZN => n58);
   U151 : INV_X1 port map( A => B(12), ZN => n57);
   U152 : NOR2_X1 port map( A1 => n59, A2 => n60, ZN => OUT_LOGIC_AND(11));
   U153 : INV_X1 port map( A => A(11), ZN => n60);
   U154 : INV_X1 port map( A => B(11), ZN => n59);
   U155 : NOR2_X1 port map( A1 => n61, A2 => n62, ZN => OUT_LOGIC_AND(10));
   U156 : INV_X1 port map( A => A(10), ZN => n62);
   U157 : INV_X1 port map( A => B(10), ZN => n61);
   U158 : NOR2_X1 port map( A1 => n63, A2 => n64, ZN => OUT_LOGIC_AND(0));
   U159 : INV_X1 port map( A => A(0), ZN => n64);
   U160 : INV_X1 port map( A => B(0), ZN => n63);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SHIFTER_GENERIC_N32 is

   port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
         downto 0);  LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE : in std_logic;  
         OUTPUT : out std_logic_vector (31 downto 0));

end SHIFTER_GENERIC_N32;

architecture SYN_BEHAVIORAL of SHIFTER_GENERIC_N32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI222_X1
      port( A1, A2, B1, B2, C1, C2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component AND3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component SHIFTER_GENERIC_N32_DW_rbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_lbsh_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_sra_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_rash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW_sla_0
      port( A : in std_logic_vector (31 downto 0);  SH : in std_logic_vector (4
            downto 0);  SH_TC : in std_logic;  B : out std_logic_vector (31 
            downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32_DW01_ash_0
      port( A : in std_logic_vector (31 downto 0);  DATA_TC : in std_logic;  SH
            : in std_logic_vector (4 downto 0);  SH_TC : in std_logic;  B : out
            std_logic_vector (31 downto 0));
   end component;
   
   signal N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, 
      N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35
      , N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49, 
      N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63, N64
      , N65, N66, N67, N68, N69, N70, N105, N106, N107, N108, N109, N110, N111,
      N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123, 
      N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134, N135, 
      N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146, N147, 
      N148, N149, N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, 
      N160, N161, N162, N163, N164, N165, N166, N167, N168, N202, N203, N204, 
      N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216, 
      N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, 
      N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240, 
      N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, 
      N253, N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264, 
      N265, n14_port, n15_port, n16_port, n17_port, n18_port, n19_port, n1, n2,
      n3, n4, n5, n6, n7_port, n8_port, n9_port, n10_port, n11_port, n12_port, 
      n13_port, n20_port, n21_port, n22_port, n23_port, n24_port, n25_port, 
      n26_port, n27_port, n28_port, n29_port, n30_port, n31_port, n32_port, 
      n33_port, n34_port, n35_port, n36_port, n37_port, n38_port, n39_port, 
      n40_port, n41_port, n42_port, n43_port, n44_port, n45_port, n46_port, 
      n47_port, n48_port, n49_port, n50_port, n51_port, n52_port, n53_port, 
      n54_port, n55_port, n56_port, n57_port, n58_port, n59_port, n60_port, 
      n61_port, n62_port, n63_port, n64_port, n65_port, n66_port, n67_port, 
      n68_port, n69_port, n70_port, n71, n72, n73, n74, n75, n76, n77, n78, n79
      : std_logic;

begin
   
   n14_port <= '0';
   n15_port <= '0';
   n16_port <= '0';
   n17_port <= '0';
   n18_port <= '0';
   n19_port <= '0';
   C88 : SHIFTER_GENERIC_N32_DW01_ash_0 port map( A(31) => A(31), A(30) => 
                           A(30), A(29) => A(29), A(28) => A(28), A(27) => 
                           A(27), A(26) => A(26), A(25) => A(25), A(24) => 
                           A(24), A(23) => A(23), A(22) => A(22), A(21) => 
                           A(21), A(20) => A(20), A(19) => A(19), A(18) => 
                           A(18), A(17) => A(17), A(16) => A(16), A(15) => 
                           A(15), A(14) => A(14), A(13) => A(13), A(12) => 
                           A(12), A(11) => A(11), A(10) => A(10), A(9) => A(9),
                           A(8) => A(8), A(7) => A(7), A(6) => A(6), A(5) => 
                           A(5), A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1)
                           => A(1), A(0) => A(0), DATA_TC => n14_port, SH(4) =>
                           n1, SH(3) => B(3), SH(2) => B(2), SH(1) => B(1), 
                           SH(0) => B(0), SH_TC => n14_port, B(31) => N265, 
                           B(30) => N264, B(29) => N263, B(28) => N262, B(27) 
                           => N261, B(26) => N260, B(25) => N259, B(24) => N258
                           , B(23) => N257, B(22) => N256, B(21) => N255, B(20)
                           => N254, B(19) => N253, B(18) => N252, B(17) => N251
                           , B(16) => N250, B(15) => N249, B(14) => N248, B(13)
                           => N247, B(12) => N246, B(11) => N245, B(10) => N244
                           , B(9) => N243, B(8) => N242, B(7) => N241, B(6) => 
                           N240, B(5) => N239, B(4) => N238, B(3) => N237, B(2)
                           => N236, B(1) => N235, B(0) => N234);
   C86 : SHIFTER_GENERIC_N32_DW_sla_0 port map( A(31) => A(31), A(30) => A(30),
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), SH(4) => n1, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n15_port, B(31) => N233, B(30) => N232, B(29) => 
                           N231, B(28) => N230, B(27) => N229, B(26) => N228, 
                           B(25) => N227, B(24) => N226, B(23) => N225, B(22) 
                           => N224, B(21) => N223, B(20) => N222, B(19) => N221
                           , B(18) => N220, B(17) => N219, B(16) => N218, B(15)
                           => N217, B(14) => N216, B(13) => N215, B(12) => N214
                           , B(11) => N213, B(10) => N212, B(9) => N211, B(8) 
                           => N210, B(7) => N209, B(6) => N208, B(5) => N207, 
                           B(4) => N206, B(3) => N205, B(2) => N204, B(1) => 
                           N203, B(0) => N202);
   C50 : SHIFTER_GENERIC_N32_DW_rash_0 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), DATA_TC => n16_port, SH(4) => n1
                           , SH(3) => B(3), SH(2) => B(2), SH(1) => B(1), SH(0)
                           => B(0), SH_TC => n16_port, B(31) => N168, B(30) => 
                           N167, B(29) => N166, B(28) => N165, B(27) => N164, 
                           B(26) => N163, B(25) => N162, B(24) => N161, B(23) 
                           => N160, B(22) => N159, B(21) => N158, B(20) => N157
                           , B(19) => N156, B(18) => N155, B(17) => N154, B(16)
                           => N153, B(15) => N152, B(14) => N151, B(13) => N150
                           , B(12) => N149, B(11) => N148, B(10) => N147, B(9) 
                           => N146, B(8) => N145, B(7) => N144, B(6) => N143, 
                           B(5) => N142, B(4) => N141, B(3) => N140, B(2) => 
                           N139, B(1) => N138, B(0) => N137);
   C48 : SHIFTER_GENERIC_N32_DW_sra_0 port map( A(31) => A(31), A(30) => A(30),
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), SH(4) => n1, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n17_port, B(31) => N136, B(30) => N135, B(29) => 
                           N134, B(28) => N133, B(27) => N132, B(26) => N131, 
                           B(25) => N130, B(24) => N129, B(23) => N128, B(22) 
                           => N127, B(21) => N126, B(20) => N125, B(19) => N124
                           , B(18) => N123, B(17) => N122, B(16) => N121, B(15)
                           => N120, B(14) => N119, B(13) => N118, B(12) => N117
                           , B(11) => N116, B(10) => N115, B(9) => N114, B(8) 
                           => N113, B(7) => N112, B(6) => N111, B(5) => N110, 
                           B(4) => N109, B(3) => N108, B(2) => N107, B(1) => 
                           N106, B(0) => N105);
   C10 : SHIFTER_GENERIC_N32_DW_lbsh_0 port map( A(31) => A(31), A(30) => A(30)
                           , A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), SH(4) => n1, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n18_port, B(31) => N70, B(30) => N69, B(29) => 
                           N68, B(28) => N67, B(27) => N66, B(26) => N65, B(25)
                           => N64, B(24) => N63, B(23) => N62, B(22) => N61, 
                           B(21) => N60, B(20) => N59, B(19) => N58, B(18) => 
                           N57, B(17) => N56, B(16) => N55, B(15) => N54, B(14)
                           => N53, B(13) => N52, B(12) => N51, B(11) => N50, 
                           B(10) => N49, B(9) => N48, B(8) => N47, B(7) => N46,
                           B(6) => N45, B(5) => N44, B(4) => N43, B(3) => N42, 
                           B(2) => N41, B(1) => N40, B(0) => N39);
   C8 : SHIFTER_GENERIC_N32_DW_rbsh_0 port map( A(31) => A(31), A(30) => A(30),
                           A(29) => A(29), A(28) => A(28), A(27) => A(27), 
                           A(26) => A(26), A(25) => A(25), A(24) => A(24), 
                           A(23) => A(23), A(22) => A(22), A(21) => A(21), 
                           A(20) => A(20), A(19) => A(19), A(18) => A(18), 
                           A(17) => A(17), A(16) => A(16), A(15) => A(15), 
                           A(14) => A(14), A(13) => A(13), A(12) => A(12), 
                           A(11) => A(11), A(10) => A(10), A(9) => A(9), A(8) 
                           => A(8), A(7) => A(7), A(6) => A(6), A(5) => A(5), 
                           A(4) => A(4), A(3) => A(3), A(2) => A(2), A(1) => 
                           A(1), A(0) => A(0), SH(4) => n1, SH(3) => B(3), 
                           SH(2) => B(2), SH(1) => B(1), SH(0) => B(0), SH_TC 
                           => n19_port, B(31) => N38, B(30) => N37, B(29) => 
                           N36, B(28) => N35, B(27) => N34, B(26) => N33, B(25)
                           => N32, B(24) => N31, B(23) => N30, B(22) => N29, 
                           B(21) => N28, B(20) => N27, B(19) => N26, B(18) => 
                           N25, B(17) => N24, B(16) => N23, B(15) => N22, B(14)
                           => N21, B(13) => N20, B(12) => N19, B(11) => N18, 
                           B(10) => N17, B(9) => N16, B(8) => N15, B(7) => N14,
                           B(6) => N13, B(5) => N12, B(4) => N11, B(3) => N10, 
                           B(2) => N9, B(1) => N8, B(0) => N7);
   U5 : NOR2_X4 port map( A1 => n78, A2 => SHIFT_ROTATE, ZN => n7_port);
   U6 : NOR2_X4 port map( A1 => LEFT_RIGHT, A2 => SHIFT_ROTATE, ZN => n8_port);
   U7 : AND3_X2 port map( A1 => n78, A2 => n79, A3 => SHIFT_ROTATE, ZN => n6);
   U8 : AND3_X2 port map( A1 => SHIFT_ROTATE, A2 => LOGIC_ARITH, A3 => 
                           LEFT_RIGHT, ZN => n9_port);
   U9 : AND3_X2 port map( A1 => LOGIC_ARITH, A2 => n78, A3 => SHIFT_ROTATE, ZN 
                           => n5);
   U10 : AND3_X2 port map( A1 => SHIFT_ROTATE, A2 => n79, A3 => LEFT_RIGHT, ZN 
                           => n4);
   U13 : CLKBUF_X3 port map( A => B(4), Z => n1);
   U14 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => OUTPUT(9));
   U15 : AOI222_X1 port map( A1 => N211, A2 => n4, B1 => N146, B2 => n5, C1 => 
                           N114, C2 => n6, ZN => n3);
   U16 : AOI222_X1 port map( A1 => N48, A2 => n7_port, B1 => N16, B2 => n8_port
                           , C1 => N243, C2 => n9_port, ZN => n2);
   U17 : NAND2_X1 port map( A1 => n10_port, A2 => n11_port, ZN => OUTPUT(8));
   U18 : AOI222_X1 port map( A1 => N210, A2 => n4, B1 => N145, B2 => n5, C1 => 
                           N113, C2 => n6, ZN => n11_port);
   U19 : AOI222_X1 port map( A1 => N47, A2 => n7_port, B1 => N15, B2 => n8_port
                           , C1 => N242, C2 => n9_port, ZN => n10_port);
   U20 : NAND2_X1 port map( A1 => n12_port, A2 => n13_port, ZN => OUTPUT(7));
   U21 : AOI222_X1 port map( A1 => N209, A2 => n4, B1 => N144, B2 => n5, C1 => 
                           N112, C2 => n6, ZN => n13_port);
   U22 : AOI222_X1 port map( A1 => N46, A2 => n7_port, B1 => N14, B2 => n8_port
                           , C1 => N241, C2 => n9_port, ZN => n12_port);
   U23 : NAND2_X1 port map( A1 => n20_port, A2 => n21_port, ZN => OUTPUT(6));
   U24 : AOI222_X1 port map( A1 => N208, A2 => n4, B1 => N143, B2 => n5, C1 => 
                           N111, C2 => n6, ZN => n21_port);
   U25 : AOI222_X1 port map( A1 => N45, A2 => n7_port, B1 => N13, B2 => n8_port
                           , C1 => N240, C2 => n9_port, ZN => n20_port);
   U26 : NAND2_X1 port map( A1 => n22_port, A2 => n23_port, ZN => OUTPUT(5));
   U27 : AOI222_X1 port map( A1 => N207, A2 => n4, B1 => N142, B2 => n5, C1 => 
                           N110, C2 => n6, ZN => n23_port);
   U28 : AOI222_X1 port map( A1 => N44, A2 => n7_port, B1 => N12, B2 => n8_port
                           , C1 => N239, C2 => n9_port, ZN => n22_port);
   U29 : NAND2_X1 port map( A1 => n24_port, A2 => n25_port, ZN => OUTPUT(4));
   U30 : AOI222_X1 port map( A1 => N206, A2 => n4, B1 => N141, B2 => n5, C1 => 
                           N109, C2 => n6, ZN => n25_port);
   U31 : AOI222_X1 port map( A1 => N43, A2 => n7_port, B1 => N11, B2 => n8_port
                           , C1 => N238, C2 => n9_port, ZN => n24_port);
   U32 : NAND2_X1 port map( A1 => n26_port, A2 => n27_port, ZN => OUTPUT(3));
   U33 : AOI222_X1 port map( A1 => N205, A2 => n4, B1 => N140, B2 => n5, C1 => 
                           N108, C2 => n6, ZN => n27_port);
   U34 : AOI222_X1 port map( A1 => N42, A2 => n7_port, B1 => N10, B2 => n8_port
                           , C1 => N237, C2 => n9_port, ZN => n26_port);
   U35 : NAND2_X1 port map( A1 => n28_port, A2 => n29_port, ZN => OUTPUT(31));
   U36 : AOI222_X1 port map( A1 => N233, A2 => n4, B1 => N168, B2 => n5, C1 => 
                           N136, C2 => n6, ZN => n29_port);
   U37 : AOI222_X1 port map( A1 => N70, A2 => n7_port, B1 => N38, B2 => n8_port
                           , C1 => N265, C2 => n9_port, ZN => n28_port);
   U38 : NAND2_X1 port map( A1 => n30_port, A2 => n31_port, ZN => OUTPUT(30));
   U39 : AOI222_X1 port map( A1 => N232, A2 => n4, B1 => N167, B2 => n5, C1 => 
                           N135, C2 => n6, ZN => n31_port);
   U40 : AOI222_X1 port map( A1 => N69, A2 => n7_port, B1 => N37, B2 => n8_port
                           , C1 => N264, C2 => n9_port, ZN => n30_port);
   U41 : NAND2_X1 port map( A1 => n32_port, A2 => n33_port, ZN => OUTPUT(2));
   U42 : AOI222_X1 port map( A1 => N204, A2 => n4, B1 => N139, B2 => n5, C1 => 
                           N107, C2 => n6, ZN => n33_port);
   U43 : AOI222_X1 port map( A1 => N41, A2 => n7_port, B1 => N9, B2 => n8_port,
                           C1 => N236, C2 => n9_port, ZN => n32_port);
   U44 : NAND2_X1 port map( A1 => n34_port, A2 => n35_port, ZN => OUTPUT(29));
   U45 : AOI222_X1 port map( A1 => N231, A2 => n4, B1 => N166, B2 => n5, C1 => 
                           N134, C2 => n6, ZN => n35_port);
   U46 : AOI222_X1 port map( A1 => N68, A2 => n7_port, B1 => N36, B2 => n8_port
                           , C1 => N263, C2 => n9_port, ZN => n34_port);
   U47 : NAND2_X1 port map( A1 => n36_port, A2 => n37_port, ZN => OUTPUT(28));
   U48 : AOI222_X1 port map( A1 => N230, A2 => n4, B1 => N165, B2 => n5, C1 => 
                           N133, C2 => n6, ZN => n37_port);
   U49 : AOI222_X1 port map( A1 => N67, A2 => n7_port, B1 => N35, B2 => n8_port
                           , C1 => N262, C2 => n9_port, ZN => n36_port);
   U50 : NAND2_X1 port map( A1 => n38_port, A2 => n39_port, ZN => OUTPUT(27));
   U51 : AOI222_X1 port map( A1 => N229, A2 => n4, B1 => N164, B2 => n5, C1 => 
                           N132, C2 => n6, ZN => n39_port);
   U52 : AOI222_X1 port map( A1 => N66, A2 => n7_port, B1 => N34, B2 => n8_port
                           , C1 => N261, C2 => n9_port, ZN => n38_port);
   U53 : NAND2_X1 port map( A1 => n40_port, A2 => n41_port, ZN => OUTPUT(26));
   U54 : AOI222_X1 port map( A1 => N228, A2 => n4, B1 => N163, B2 => n5, C1 => 
                           N131, C2 => n6, ZN => n41_port);
   U55 : AOI222_X1 port map( A1 => N65, A2 => n7_port, B1 => N33, B2 => n8_port
                           , C1 => N260, C2 => n9_port, ZN => n40_port);
   U56 : NAND2_X1 port map( A1 => n42_port, A2 => n43_port, ZN => OUTPUT(25));
   U57 : AOI222_X1 port map( A1 => N227, A2 => n4, B1 => N162, B2 => n5, C1 => 
                           N130, C2 => n6, ZN => n43_port);
   U58 : AOI222_X1 port map( A1 => N64, A2 => n7_port, B1 => N32, B2 => n8_port
                           , C1 => N259, C2 => n9_port, ZN => n42_port);
   U59 : NAND2_X1 port map( A1 => n44_port, A2 => n45_port, ZN => OUTPUT(24));
   U60 : AOI222_X1 port map( A1 => N226, A2 => n4, B1 => N161, B2 => n5, C1 => 
                           N129, C2 => n6, ZN => n45_port);
   U61 : AOI222_X1 port map( A1 => N63, A2 => n7_port, B1 => N31, B2 => n8_port
                           , C1 => N258, C2 => n9_port, ZN => n44_port);
   U62 : NAND2_X1 port map( A1 => n46_port, A2 => n47_port, ZN => OUTPUT(23));
   U63 : AOI222_X1 port map( A1 => N225, A2 => n4, B1 => N160, B2 => n5, C1 => 
                           N128, C2 => n6, ZN => n47_port);
   U64 : AOI222_X1 port map( A1 => N62, A2 => n7_port, B1 => N30, B2 => n8_port
                           , C1 => N257, C2 => n9_port, ZN => n46_port);
   U65 : NAND2_X1 port map( A1 => n48_port, A2 => n49_port, ZN => OUTPUT(22));
   U66 : AOI222_X1 port map( A1 => N224, A2 => n4, B1 => N159, B2 => n5, C1 => 
                           N127, C2 => n6, ZN => n49_port);
   U67 : AOI222_X1 port map( A1 => N61, A2 => n7_port, B1 => N29, B2 => n8_port
                           , C1 => N256, C2 => n9_port, ZN => n48_port);
   U68 : NAND2_X1 port map( A1 => n50_port, A2 => n51_port, ZN => OUTPUT(21));
   U69 : AOI222_X1 port map( A1 => N223, A2 => n4, B1 => N158, B2 => n5, C1 => 
                           N126, C2 => n6, ZN => n51_port);
   U70 : AOI222_X1 port map( A1 => N60, A2 => n7_port, B1 => N28, B2 => n8_port
                           , C1 => N255, C2 => n9_port, ZN => n50_port);
   U71 : NAND2_X1 port map( A1 => n52_port, A2 => n53_port, ZN => OUTPUT(20));
   U72 : AOI222_X1 port map( A1 => N222, A2 => n4, B1 => N157, B2 => n5, C1 => 
                           N125, C2 => n6, ZN => n53_port);
   U73 : AOI222_X1 port map( A1 => N59, A2 => n7_port, B1 => N27, B2 => n8_port
                           , C1 => N254, C2 => n9_port, ZN => n52_port);
   U74 : NAND2_X1 port map( A1 => n54_port, A2 => n55_port, ZN => OUTPUT(1));
   U75 : AOI222_X1 port map( A1 => N203, A2 => n4, B1 => N138, B2 => n5, C1 => 
                           N106, C2 => n6, ZN => n55_port);
   U76 : AOI222_X1 port map( A1 => N40, A2 => n7_port, B1 => N8, B2 => n8_port,
                           C1 => N235, C2 => n9_port, ZN => n54_port);
   U77 : NAND2_X1 port map( A1 => n56_port, A2 => n57_port, ZN => OUTPUT(19));
   U78 : AOI222_X1 port map( A1 => N221, A2 => n4, B1 => N156, B2 => n5, C1 => 
                           N124, C2 => n6, ZN => n57_port);
   U79 : AOI222_X1 port map( A1 => N58, A2 => n7_port, B1 => N26, B2 => n8_port
                           , C1 => N253, C2 => n9_port, ZN => n56_port);
   U80 : NAND2_X1 port map( A1 => n58_port, A2 => n59_port, ZN => OUTPUT(18));
   U81 : AOI222_X1 port map( A1 => N220, A2 => n4, B1 => N155, B2 => n5, C1 => 
                           N123, C2 => n6, ZN => n59_port);
   U82 : AOI222_X1 port map( A1 => N57, A2 => n7_port, B1 => N25, B2 => n8_port
                           , C1 => N252, C2 => n9_port, ZN => n58_port);
   U83 : NAND2_X1 port map( A1 => n60_port, A2 => n61_port, ZN => OUTPUT(17));
   U84 : AOI222_X1 port map( A1 => N219, A2 => n4, B1 => N154, B2 => n5, C1 => 
                           N122, C2 => n6, ZN => n61_port);
   U85 : AOI222_X1 port map( A1 => N56, A2 => n7_port, B1 => N24, B2 => n8_port
                           , C1 => N251, C2 => n9_port, ZN => n60_port);
   U86 : NAND2_X1 port map( A1 => n62_port, A2 => n63_port, ZN => OUTPUT(16));
   U87 : AOI222_X1 port map( A1 => N218, A2 => n4, B1 => N153, B2 => n5, C1 => 
                           N121, C2 => n6, ZN => n63_port);
   U88 : AOI222_X1 port map( A1 => N55, A2 => n7_port, B1 => N23, B2 => n8_port
                           , C1 => N250, C2 => n9_port, ZN => n62_port);
   U89 : NAND2_X1 port map( A1 => n64_port, A2 => n65_port, ZN => OUTPUT(15));
   U90 : AOI222_X1 port map( A1 => N217, A2 => n4, B1 => N152, B2 => n5, C1 => 
                           N120, C2 => n6, ZN => n65_port);
   U91 : AOI222_X1 port map( A1 => N54, A2 => n7_port, B1 => N22, B2 => n8_port
                           , C1 => N249, C2 => n9_port, ZN => n64_port);
   U92 : NAND2_X1 port map( A1 => n66_port, A2 => n67_port, ZN => OUTPUT(14));
   U93 : AOI222_X1 port map( A1 => N216, A2 => n4, B1 => N151, B2 => n5, C1 => 
                           N119, C2 => n6, ZN => n67_port);
   U94 : AOI222_X1 port map( A1 => N53, A2 => n7_port, B1 => N21, B2 => n8_port
                           , C1 => N248, C2 => n9_port, ZN => n66_port);
   U95 : NAND2_X1 port map( A1 => n68_port, A2 => n69_port, ZN => OUTPUT(13));
   U96 : AOI222_X1 port map( A1 => N215, A2 => n4, B1 => N150, B2 => n5, C1 => 
                           N118, C2 => n6, ZN => n69_port);
   U97 : AOI222_X1 port map( A1 => N52, A2 => n7_port, B1 => N20, B2 => n8_port
                           , C1 => N247, C2 => n9_port, ZN => n68_port);
   U98 : NAND2_X1 port map( A1 => n70_port, A2 => n71, ZN => OUTPUT(12));
   U99 : AOI222_X1 port map( A1 => N214, A2 => n4, B1 => N149, B2 => n5, C1 => 
                           N117, C2 => n6, ZN => n71);
   U100 : AOI222_X1 port map( A1 => N51, A2 => n7_port, B1 => N19, B2 => 
                           n8_port, C1 => N246, C2 => n9_port, ZN => n70_port);
   U101 : NAND2_X1 port map( A1 => n72, A2 => n73, ZN => OUTPUT(11));
   U102 : AOI222_X1 port map( A1 => N213, A2 => n4, B1 => N148, B2 => n5, C1 =>
                           N116, C2 => n6, ZN => n73);
   U103 : AOI222_X1 port map( A1 => N50, A2 => n7_port, B1 => N18, B2 => 
                           n8_port, C1 => N245, C2 => n9_port, ZN => n72);
   U104 : NAND2_X1 port map( A1 => n74, A2 => n75, ZN => OUTPUT(10));
   U105 : AOI222_X1 port map( A1 => N212, A2 => n4, B1 => N147, B2 => n5, C1 =>
                           N115, C2 => n6, ZN => n75);
   U106 : AOI222_X1 port map( A1 => N49, A2 => n7_port, B1 => N17, B2 => 
                           n8_port, C1 => N244, C2 => n9_port, ZN => n74);
   U107 : NAND2_X1 port map( A1 => n76, A2 => n77, ZN => OUTPUT(0));
   U108 : AOI222_X1 port map( A1 => N202, A2 => n4, B1 => N137, B2 => n5, C1 =>
                           N105, C2 => n6, ZN => n77);
   U109 : INV_X1 port map( A => LOGIC_ARITH, ZN => n79);
   U110 : AOI222_X1 port map( A1 => N39, A2 => n7_port, B1 => N7, B2 => n8_port
                           , C1 => N234, C2 => n9_port, ZN => n76);
   U111 : INV_X1 port map( A => LEFT_RIGHT, ZN => n78);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity RCA_GEN_NBIT32 is

   port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (31 downto 0);  Co : out std_logic);

end RCA_GEN_NBIT32;

architecture SYN_structural of RCA_GEN_NBIT32 is

   component FA_65
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_66
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_67
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_68
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_69
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_70
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_71
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_72
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_73
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_74
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_75
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_76
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_77
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_78
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_79
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_80
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_81
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_82
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_83
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_84
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_85
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_86
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_87
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_88
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_89
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_90
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_91
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_92
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_93
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_94
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_95
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal CTMP_31_port, CTMP_30_port, CTMP_29_port, CTMP_28_port, CTMP_27_port,
      CTMP_26_port, CTMP_25_port, CTMP_24_port, CTMP_23_port, CTMP_22_port, 
      CTMP_21_port, CTMP_20_port, CTMP_19_port, CTMP_18_port, CTMP_17_port, 
      CTMP_16_port, CTMP_15_port, CTMP_14_port, CTMP_13_port, CTMP_12_port, 
      CTMP_11_port, CTMP_10_port, CTMP_9_port, CTMP_8_port, CTMP_7_port, 
      CTMP_6_port, CTMP_5_port, CTMP_4_port, CTMP_3_port, CTMP_2_port, 
      CTMP_1_port : std_logic;

begin
   
   fai_1 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           CTMP_1_port);
   fai_2 : FA_95 port map( A => A(1), B => B(1), Ci => CTMP_1_port, S => S(1), 
                           Co => CTMP_2_port);
   fai_3 : FA_94 port map( A => A(2), B => B(2), Ci => CTMP_2_port, S => S(2), 
                           Co => CTMP_3_port);
   fai_4 : FA_93 port map( A => A(3), B => B(3), Ci => CTMP_3_port, S => S(3), 
                           Co => CTMP_4_port);
   fai_5 : FA_92 port map( A => A(4), B => B(4), Ci => CTMP_4_port, S => S(4), 
                           Co => CTMP_5_port);
   fai_6 : FA_91 port map( A => A(5), B => B(5), Ci => CTMP_5_port, S => S(5), 
                           Co => CTMP_6_port);
   fai_7 : FA_90 port map( A => A(6), B => B(6), Ci => CTMP_6_port, S => S(6), 
                           Co => CTMP_7_port);
   fai_8 : FA_89 port map( A => A(7), B => B(7), Ci => CTMP_7_port, S => S(7), 
                           Co => CTMP_8_port);
   fai_9 : FA_88 port map( A => A(8), B => B(8), Ci => CTMP_8_port, S => S(8), 
                           Co => CTMP_9_port);
   fai_10 : FA_87 port map( A => A(9), B => B(9), Ci => CTMP_9_port, S => S(9),
                           Co => CTMP_10_port);
   fai_11 : FA_86 port map( A => A(10), B => B(10), Ci => CTMP_10_port, S => 
                           S(10), Co => CTMP_11_port);
   fai_12 : FA_85 port map( A => A(11), B => B(11), Ci => CTMP_11_port, S => 
                           S(11), Co => CTMP_12_port);
   fai_13 : FA_84 port map( A => A(12), B => B(12), Ci => CTMP_12_port, S => 
                           S(12), Co => CTMP_13_port);
   fai_14 : FA_83 port map( A => A(13), B => B(13), Ci => CTMP_13_port, S => 
                           S(13), Co => CTMP_14_port);
   fai_15 : FA_82 port map( A => A(14), B => B(14), Ci => CTMP_14_port, S => 
                           S(14), Co => CTMP_15_port);
   fai_16 : FA_81 port map( A => A(15), B => B(15), Ci => CTMP_15_port, S => 
                           S(15), Co => CTMP_16_port);
   fai_17 : FA_80 port map( A => A(16), B => B(16), Ci => CTMP_16_port, S => 
                           S(16), Co => CTMP_17_port);
   fai_18 : FA_79 port map( A => A(17), B => B(17), Ci => CTMP_17_port, S => 
                           S(17), Co => CTMP_18_port);
   fai_19 : FA_78 port map( A => A(18), B => B(18), Ci => CTMP_18_port, S => 
                           S(18), Co => CTMP_19_port);
   fai_20 : FA_77 port map( A => A(19), B => B(19), Ci => CTMP_19_port, S => 
                           S(19), Co => CTMP_20_port);
   fai_21 : FA_76 port map( A => A(20), B => B(20), Ci => CTMP_20_port, S => 
                           S(20), Co => CTMP_21_port);
   fai_22 : FA_75 port map( A => A(21), B => B(21), Ci => CTMP_21_port, S => 
                           S(21), Co => CTMP_22_port);
   fai_23 : FA_74 port map( A => A(22), B => B(22), Ci => CTMP_22_port, S => 
                           S(22), Co => CTMP_23_port);
   fai_24 : FA_73 port map( A => A(23), B => B(23), Ci => CTMP_23_port, S => 
                           S(23), Co => CTMP_24_port);
   fai_25 : FA_72 port map( A => A(24), B => B(24), Ci => CTMP_24_port, S => 
                           S(24), Co => CTMP_25_port);
   fai_26 : FA_71 port map( A => A(25), B => B(25), Ci => CTMP_25_port, S => 
                           S(25), Co => CTMP_26_port);
   fai_27 : FA_70 port map( A => A(26), B => B(26), Ci => CTMP_26_port, S => 
                           S(26), Co => CTMP_27_port);
   fai_28 : FA_69 port map( A => A(27), B => B(27), Ci => CTMP_27_port, S => 
                           S(27), Co => CTMP_28_port);
   fai_29 : FA_68 port map( A => A(28), B => B(28), Ci => CTMP_28_port, S => 
                           S(28), Co => CTMP_29_port);
   fai_30 : FA_67 port map( A => A(29), B => B(29), Ci => CTMP_29_port, S => 
                           S(29), Co => CTMP_30_port);
   fai_31 : FA_66 port map( A => A(30), B => B(30), Ci => CTMP_30_port, S => 
                           S(30), Co => CTMP_31_port);
   fai_32 : FA_65 port map( A => A(31), B => B(31), Ci => CTMP_31_port, S => 
                           S(31), Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_N5 is

   port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : out
         std_logic_vector (4 downto 0));

end mux21_N5;

architecture SYN_behavioural of mux21_N5 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U2 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U3 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U4 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U5 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity AluOpCodeGen is

   port( IR_opcode : in std_logic_vector (5 downto 0);  IR_func : in 
         std_logic_vector (10 downto 0);  AluOpCode : out std_logic_vector (2 
         downto 0);  Add_Subn : out std_logic;  CompareCode : out 
         std_logic_vector (3 downto 0);  ShiftOpCode : out std_logic_vector (2 
         downto 0));

end AluOpCodeGen;

architecture SYN_beh of AluOpCodeGen is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI33_X1
      port( A1, A2, A3, B1, B2, B3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X2
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   signal n37, ShiftOpCode_0_port, ShiftOpCode_1_port, n2, n3, n4, n5, n6, n7, 
      n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, 
      n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36 : 
      std_logic;

begin
   ShiftOpCode <= ( ShiftOpCode_0_port, ShiftOpCode_1_port, ShiftOpCode_0_port 
      );
   
   U3 : CLKBUF_X2 port map( A => n37, Z => Add_Subn);
   U4 : OAI22_X1 port map( A1 => IR_func(1), A2 => n2, B1 => IR_opcode(1), B2 
                           => n3, ZN => ShiftOpCode_1_port);
   U5 : NOR3_X1 port map( A1 => n4, A2 => IR_opcode(3), A3 => IR_opcode(0), ZN 
                           => CompareCode(3));
   U6 : NOR3_X1 port map( A1 => n5, A2 => IR_opcode(3), A3 => n4, ZN => 
                           CompareCode(2));
   U7 : OAI21_X1 port map( B1 => n6, B2 => n7, A => n8, ZN => CompareCode(1));
   U8 : OR3_X1 port map( A1 => n9, A2 => n10, A3 => n11, ZN => n8);
   U9 : OAI21_X1 port map( B1 => IR_func(2), B2 => n7, A => n12, ZN => 
                           CompareCode(0));
   U10 : NAND3_X1 port map( A1 => IR_opcode(4), A2 => n10, A3 => n13, ZN => n12
                           );
   U11 : OAI211_X1 port map( C1 => n14, C2 => n11, A => n7, B => n15, ZN => 
                           AluOpCode(2));
   U12 : NAND2_X1 port map( A1 => IR_func(3), A2 => n16, ZN => n7);
   U13 : INV_X1 port map( A => n17, ZN => n16);
   U14 : INV_X1 port map( A => n13, ZN => n11);
   U15 : NOR4_X1 port map( A1 => n18, A2 => n5, A3 => IR_opcode(1), A4 => 
                           IR_opcode(5), ZN => n13);
   U16 : INV_X1 port map( A => n19, ZN => AluOpCode(1));
   U17 : AOI21_X1 port map( B1 => n20, B2 => IR_func(2), A => n9, ZN => n19);
   U18 : OAI33_X1 port map( A1 => n18, A2 => n4, A3 => n5, B1 => n21, B2 => n10
                           , B3 => n22, ZN => n9);
   U19 : OAI22_X1 port map( A1 => n17, A2 => IR_func(3), B1 => n23, B2 => n24, 
                           ZN => n20);
   U20 : NAND4_X1 port map( A1 => IR_func(5), A2 => IR_func(0), A3 => n25, A4 
                           => n23, ZN => n17);
   U21 : OAI221_X1 port map( B1 => n26, B2 => n22, C1 => n6, C2 => n24, A => 
                           n15, ZN => AluOpCode(0));
   U22 : INV_X1 port map( A => ShiftOpCode_0_port, ZN => n15);
   U23 : NAND2_X1 port map( A1 => n2, A2 => n3, ZN => ShiftOpCode_0_port);
   U24 : NAND4_X1 port map( A1 => IR_opcode(4), A2 => IR_opcode(2), A3 => n27, 
                           A4 => n5, ZN => n3);
   U25 : NOR2_X1 port map( A1 => IR_opcode(5), A2 => IR_opcode(3), ZN => n27);
   U26 : NAND3_X1 port map( A1 => n28, A2 => n29, A3 => IR_func(2), ZN => n2);
   U27 : INV_X1 port map( A => IR_func(5), ZN => n29);
   U28 : INV_X1 port map( A => IR_func(2), ZN => n6);
   U29 : INV_X1 port map( A => n30, ZN => n26);
   U30 : OAI21_X1 port map( B1 => n21, B2 => n10, A => n4, ZN => n30);
   U31 : OR2_X1 port map( A1 => n31, A2 => n10, ZN => n4);
   U32 : OAI33_X1 port map( A1 => n23, A2 => IR_func(2), A3 => n24, B1 => n21, 
                           B2 => IR_opcode(2), B3 => n22, ZN => n37);
   U33 : NAND2_X1 port map( A1 => IR_opcode(3), A2 => n5, ZN => n22);
   U34 : NAND3_X1 port map( A1 => n14, A2 => n32, A3 => IR_opcode(1), ZN => n21
                           );
   U35 : INV_X1 port map( A => IR_opcode(5), ZN => n32);
   U36 : INV_X1 port map( A => IR_opcode(4), ZN => n14);
   U37 : NAND2_X1 port map( A1 => IR_func(5), A2 => n28, ZN => n24);
   U38 : NOR3_X1 port map( A1 => IR_func(0), A2 => IR_func(3), A3 => n33, ZN =>
                           n28);
   U39 : INV_X1 port map( A => n25, ZN => n33);
   U40 : NOR4_X1 port map( A1 => IR_func(10), A2 => n31, A3 => n34, A4 => n35, 
                           ZN => n25);
   U41 : NAND4_X1 port map( A1 => n10, A2 => n18, A3 => n5, A4 => n36, ZN => 
                           n35);
   U42 : NOR2_X1 port map( A1 => IR_func(9), A2 => IR_func(8), ZN => n36);
   U43 : INV_X1 port map( A => IR_opcode(0), ZN => n5);
   U44 : INV_X1 port map( A => IR_opcode(3), ZN => n18);
   U45 : INV_X1 port map( A => IR_opcode(2), ZN => n10);
   U46 : OR3_X1 port map( A1 => IR_func(7), A2 => IR_func(6), A3 => IR_func(4),
                           ZN => n34);
   U47 : OR3_X1 port map( A1 => IR_opcode(4), A2 => IR_opcode(5), A3 => 
                           IR_opcode(1), ZN => n31);
   U48 : INV_X1 port map( A => IR_func(1), ZN => n23);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity ALU_N32 is

   port( AluOpCode : in std_logic_vector (2 downto 0);  CompareOpCode : in 
         std_logic_vector (3 downto 0);  Add_subn : in std_logic;  ShiftOpCode 
         : in std_logic_vector (2 downto 0);  DATA1, DATA2 : in 
         std_logic_vector (31 downto 0);  OUTALU, return_address : out 
         std_logic_vector (31 downto 0);  CompBranch : out std_logic);

end ALU_N32;

architecture SYN_BEHAVIOR of ALU_N32 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX_6to1_n32
      port( A, B, C, D, E, F : in std_logic_vector (31 downto 0);  S : in 
            std_logic_vector (2 downto 0);  Y : out std_logic_vector (31 downto
            0));
   end component;
   
   component MUX_2to1_n32
      port( A, B : in std_logic_vector (31 downto 0);  S : in std_logic;  Y : 
            out std_logic_vector (31 downto 0));
   end component;
   
   component compare_N32
      port( num1, num2 : in std_logic_vector (31 downto 0);  less, equal, 
            greater : out std_logic);
   end component;
   
   component p4_adder_N32_N_carry4
      port( A, B : in std_logic_vector (31 downto 0);  Cin : in std_logic;  SUM
            : out std_logic_vector (31 downto 0));
   end component;
   
   component operatore_logic_REG_SIZE32
      port( A, B : in std_logic_vector (31 downto 0);  OUT_LOGIC_AND, 
            OUT_LOGIC_OR, OUT_LOGIC_XOR : out std_logic_vector (31 downto 0));
   end component;
   
   component SHIFTER_GENERIC_N32
      port( A : in std_logic_vector (31 downto 0);  B : in std_logic_vector (4 
            downto 0);  LOGIC_ARITH, LEFT_RIGHT, SHIFT_ROTATE : in std_logic;  
            OUTPUT : out std_logic_vector (31 downto 0));
   end component;
   
   component RCA_GEN_NBIT32
      port( A, B : in std_logic_vector (31 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (31 downto 0);  Co : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, shift_out_31_port, shift_out_30_port, 
      shift_out_29_port, shift_out_28_port, shift_out_27_port, 
      shift_out_26_port, shift_out_25_port, shift_out_24_port, 
      shift_out_23_port, shift_out_22_port, shift_out_21_port, 
      shift_out_20_port, shift_out_19_port, shift_out_18_port, 
      shift_out_17_port, shift_out_16_port, shift_out_15_port, 
      shift_out_14_port, shift_out_13_port, shift_out_12_port, 
      shift_out_11_port, shift_out_10_port, shift_out_9_port, shift_out_8_port,
      shift_out_7_port, shift_out_6_port, shift_out_5_port, shift_out_4_port, 
      shift_out_3_port, shift_out_2_port, shift_out_1_port, shift_out_0_port, 
      AND_OUT_31_port, AND_OUT_30_port, AND_OUT_29_port, AND_OUT_28_port, 
      AND_OUT_27_port, AND_OUT_26_port, AND_OUT_25_port, AND_OUT_24_port, 
      AND_OUT_23_port, AND_OUT_22_port, AND_OUT_21_port, AND_OUT_20_port, 
      AND_OUT_19_port, AND_OUT_18_port, AND_OUT_17_port, AND_OUT_16_port, 
      AND_OUT_15_port, AND_OUT_14_port, AND_OUT_13_port, AND_OUT_12_port, 
      AND_OUT_11_port, AND_OUT_10_port, AND_OUT_9_port, AND_OUT_8_port, 
      AND_OUT_7_port, AND_OUT_6_port, AND_OUT_5_port, AND_OUT_4_port, 
      AND_OUT_3_port, AND_OUT_2_port, AND_OUT_1_port, AND_OUT_0_port, 
      OR_OUT_31_port, OR_OUT_30_port, OR_OUT_29_port, OR_OUT_28_port, 
      OR_OUT_27_port, OR_OUT_26_port, OR_OUT_25_port, OR_OUT_24_port, 
      OR_OUT_23_port, OR_OUT_22_port, OR_OUT_21_port, OR_OUT_20_port, 
      OR_OUT_19_port, OR_OUT_18_port, OR_OUT_17_port, OR_OUT_16_port, 
      OR_OUT_15_port, OR_OUT_14_port, OR_OUT_13_port, OR_OUT_12_port, 
      OR_OUT_11_port, OR_OUT_10_port, OR_OUT_9_port, OR_OUT_8_port, 
      OR_OUT_7_port, OR_OUT_6_port, OR_OUT_5_port, OR_OUT_4_port, OR_OUT_3_port
      , OR_OUT_2_port, OR_OUT_1_port, OR_OUT_0_port, XOR_OUT_31_port, 
      XOR_OUT_30_port, XOR_OUT_29_port, XOR_OUT_28_port, XOR_OUT_27_port, 
      XOR_OUT_26_port, XOR_OUT_25_port, XOR_OUT_24_port, XOR_OUT_23_port, 
      XOR_OUT_22_port, XOR_OUT_21_port, XOR_OUT_20_port, XOR_OUT_19_port, 
      XOR_OUT_18_port, XOR_OUT_17_port, XOR_OUT_16_port, XOR_OUT_15_port, 
      XOR_OUT_14_port, XOR_OUT_13_port, XOR_OUT_12_port, XOR_OUT_11_port, 
      XOR_OUT_10_port, XOR_OUT_9_port, XOR_OUT_8_port, XOR_OUT_7_port, 
      XOR_OUT_6_port, XOR_OUT_5_port, XOR_OUT_4_port, XOR_OUT_3_port, 
      XOR_OUT_2_port, XOR_OUT_1_port, XOR_OUT_0_port, add_sub_out_31_port, 
      add_sub_out_30_port, add_sub_out_29_port, add_sub_out_28_port, 
      add_sub_out_27_port, add_sub_out_26_port, add_sub_out_25_port, 
      add_sub_out_24_port, add_sub_out_23_port, add_sub_out_22_port, 
      add_sub_out_21_port, add_sub_out_20_port, add_sub_out_19_port, 
      add_sub_out_18_port, add_sub_out_17_port, add_sub_out_16_port, 
      add_sub_out_15_port, add_sub_out_14_port, add_sub_out_13_port, 
      add_sub_out_12_port, add_sub_out_11_port, add_sub_out_10_port, 
      add_sub_out_9_port, add_sub_out_8_port, add_sub_out_7_port, 
      add_sub_out_6_port, add_sub_out_5_port, add_sub_out_4_port, 
      add_sub_out_3_port, add_sub_out_2_port, add_sub_out_1_port, 
      add_sub_out_0_port, comp_eq, comp_greater, sel_mux_comp_out, 
      comp_out_31_port, comp_out_30_port, comp_out_29_port, comp_out_28_port, 
      comp_out_27_port, comp_out_26_port, comp_out_25_port, comp_out_24_port, 
      comp_out_23_port, comp_out_22_port, comp_out_21_port, comp_out_20_port, 
      comp_out_19_port, comp_out_18_port, comp_out_17_port, comp_out_16_port, 
      comp_out_15_port, comp_out_14_port, comp_out_13_port, comp_out_12_port, 
      comp_out_11_port, comp_out_10_port, comp_out_9_port, comp_out_8_port, 
      comp_out_7_port, comp_out_6_port, comp_out_5_port, comp_out_4_port, 
      comp_out_3_port, comp_out_2_port, comp_out_1_port, comp_out_0_port, 
      net2103, net2104, n1, n2, n3 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   adder4 : RCA_GEN_NBIT32 port map( A(31) => DATA1(31), A(30) => DATA1(30), 
                           A(29) => DATA1(29), A(28) => DATA1(28), A(27) => 
                           DATA1(27), A(26) => DATA1(26), A(25) => DATA1(25), 
                           A(24) => DATA1(24), A(23) => DATA1(23), A(22) => 
                           DATA1(22), A(21) => DATA1(21), A(20) => DATA1(20), 
                           A(19) => DATA1(19), A(18) => DATA1(18), A(17) => 
                           DATA1(17), A(16) => DATA1(16), A(15) => DATA1(15), 
                           A(14) => DATA1(14), A(13) => DATA1(13), A(12) => 
                           DATA1(12), A(11) => DATA1(11), A(10) => DATA1(10), 
                           A(9) => DATA1(9), A(8) => DATA1(8), A(7) => DATA1(7)
                           , A(6) => DATA1(6), A(5) => DATA1(5), A(4) => 
                           DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2), A(1) 
                           => DATA1(1), A(0) => DATA1(0), B(31) => 
                           X_Logic0_port, B(30) => X_Logic0_port, B(29) => 
                           X_Logic0_port, B(28) => X_Logic0_port, B(27) => 
                           X_Logic0_port, B(26) => X_Logic0_port, B(25) => 
                           X_Logic0_port, B(24) => X_Logic0_port, B(23) => 
                           X_Logic0_port, B(22) => X_Logic0_port, B(21) => 
                           X_Logic0_port, B(20) => X_Logic0_port, B(19) => 
                           X_Logic0_port, B(18) => X_Logic0_port, B(17) => 
                           X_Logic0_port, B(16) => X_Logic0_port, B(15) => 
                           X_Logic0_port, B(14) => X_Logic0_port, B(13) => 
                           X_Logic0_port, B(12) => X_Logic0_port, B(11) => 
                           X_Logic0_port, B(10) => X_Logic0_port, B(9) => 
                           X_Logic0_port, B(8) => X_Logic0_port, B(7) => 
                           X_Logic0_port, B(6) => X_Logic0_port, B(5) => 
                           X_Logic0_port, B(4) => X_Logic0_port, B(3) => 
                           X_Logic0_port, B(2) => X_Logic1_port, B(1) => 
                           X_Logic0_port, B(0) => X_Logic0_port, Ci => 
                           X_Logic0_port, S(31) => return_address(31), S(30) =>
                           return_address(30), S(29) => return_address(29), 
                           S(28) => return_address(28), S(27) => 
                           return_address(27), S(26) => return_address(26), 
                           S(25) => return_address(25), S(24) => 
                           return_address(24), S(23) => return_address(23), 
                           S(22) => return_address(22), S(21) => 
                           return_address(21), S(20) => return_address(20), 
                           S(19) => return_address(19), S(18) => 
                           return_address(18), S(17) => return_address(17), 
                           S(16) => return_address(16), S(15) => 
                           return_address(15), S(14) => return_address(14), 
                           S(13) => return_address(13), S(12) => 
                           return_address(12), S(11) => return_address(11), 
                           S(10) => return_address(10), S(9) => 
                           return_address(9), S(8) => return_address(8), S(7) 
                           => return_address(7), S(6) => return_address(6), 
                           S(5) => return_address(5), S(4) => return_address(4)
                           , S(3) => return_address(3), S(2) => 
                           return_address(2), S(1) => return_address(1), S(0) 
                           => return_address(0), Co => net2104);
   shifter : SHIFTER_GENERIC_N32 port map( A(31) => DATA1(31), A(30) => 
                           DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28), 
                           A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), B(4) => 
                           DATA2(4), B(3) => DATA2(3), B(2) => DATA2(2), B(1) 
                           => DATA2(1), B(0) => DATA2(0), LOGIC_ARITH => 
                           ShiftOpCode(2), LEFT_RIGHT => ShiftOpCode(1), 
                           SHIFT_ROTATE => ShiftOpCode(0), OUTPUT(31) => 
                           shift_out_31_port, OUTPUT(30) => shift_out_30_port, 
                           OUTPUT(29) => shift_out_29_port, OUTPUT(28) => 
                           shift_out_28_port, OUTPUT(27) => shift_out_27_port, 
                           OUTPUT(26) => shift_out_26_port, OUTPUT(25) => 
                           shift_out_25_port, OUTPUT(24) => shift_out_24_port, 
                           OUTPUT(23) => shift_out_23_port, OUTPUT(22) => 
                           shift_out_22_port, OUTPUT(21) => shift_out_21_port, 
                           OUTPUT(20) => shift_out_20_port, OUTPUT(19) => 
                           shift_out_19_port, OUTPUT(18) => shift_out_18_port, 
                           OUTPUT(17) => shift_out_17_port, OUTPUT(16) => 
                           shift_out_16_port, OUTPUT(15) => shift_out_15_port, 
                           OUTPUT(14) => shift_out_14_port, OUTPUT(13) => 
                           shift_out_13_port, OUTPUT(12) => shift_out_12_port, 
                           OUTPUT(11) => shift_out_11_port, OUTPUT(10) => 
                           shift_out_10_port, OUTPUT(9) => shift_out_9_port, 
                           OUTPUT(8) => shift_out_8_port, OUTPUT(7) => 
                           shift_out_7_port, OUTPUT(6) => shift_out_6_port, 
                           OUTPUT(5) => shift_out_5_port, OUTPUT(4) => 
                           shift_out_4_port, OUTPUT(3) => shift_out_3_port, 
                           OUTPUT(2) => shift_out_2_port, OUTPUT(1) => 
                           shift_out_1_port, OUTPUT(0) => shift_out_0_port);
   logic_operations : operatore_logic_REG_SIZE32 port map( A(31) => DATA1(31), 
                           A(30) => DATA1(30), A(29) => DATA1(29), A(28) => 
                           DATA1(28), A(27) => DATA1(27), A(26) => DATA1(26), 
                           A(25) => DATA1(25), A(24) => DATA1(24), A(23) => 
                           DATA1(23), A(22) => DATA1(22), A(21) => DATA1(21), 
                           A(20) => DATA1(20), A(19) => DATA1(19), A(18) => 
                           DATA1(18), A(17) => DATA1(17), A(16) => DATA1(16), 
                           A(15) => DATA1(15), A(14) => DATA1(14), A(13) => 
                           DATA1(13), A(12) => DATA1(12), A(11) => DATA1(11), 
                           A(10) => DATA1(10), A(9) => DATA1(9), A(8) => 
                           DATA1(8), A(7) => DATA1(7), A(6) => DATA1(6), A(5) 
                           => DATA1(5), A(4) => DATA1(4), A(3) => DATA1(3), 
                           A(2) => DATA1(2), A(1) => DATA1(1), A(0) => DATA1(0)
                           , B(31) => DATA2(31), B(30) => DATA2(30), B(29) => 
                           DATA2(29), B(28) => DATA2(28), B(27) => DATA2(27), 
                           B(26) => DATA2(26), B(25) => DATA2(25), B(24) => 
                           DATA2(24), B(23) => DATA2(23), B(22) => DATA2(22), 
                           B(21) => DATA2(21), B(20) => DATA2(20), B(19) => 
                           DATA2(19), B(18) => DATA2(18), B(17) => DATA2(17), 
                           B(16) => DATA2(16), B(15) => DATA2(15), B(14) => 
                           DATA2(14), B(13) => DATA2(13), B(12) => DATA2(12), 
                           B(11) => DATA2(11), B(10) => DATA2(10), B(9) => 
                           DATA2(9), B(8) => DATA2(8), B(7) => DATA2(7), B(6) 
                           => DATA2(6), B(5) => DATA2(5), B(4) => DATA2(4), 
                           B(3) => DATA2(3), B(2) => DATA2(2), B(1) => DATA2(1)
                           , B(0) => DATA2(0), OUT_LOGIC_AND(31) => 
                           AND_OUT_31_port, OUT_LOGIC_AND(30) => 
                           AND_OUT_30_port, OUT_LOGIC_AND(29) => 
                           AND_OUT_29_port, OUT_LOGIC_AND(28) => 
                           AND_OUT_28_port, OUT_LOGIC_AND(27) => 
                           AND_OUT_27_port, OUT_LOGIC_AND(26) => 
                           AND_OUT_26_port, OUT_LOGIC_AND(25) => 
                           AND_OUT_25_port, OUT_LOGIC_AND(24) => 
                           AND_OUT_24_port, OUT_LOGIC_AND(23) => 
                           AND_OUT_23_port, OUT_LOGIC_AND(22) => 
                           AND_OUT_22_port, OUT_LOGIC_AND(21) => 
                           AND_OUT_21_port, OUT_LOGIC_AND(20) => 
                           AND_OUT_20_port, OUT_LOGIC_AND(19) => 
                           AND_OUT_19_port, OUT_LOGIC_AND(18) => 
                           AND_OUT_18_port, OUT_LOGIC_AND(17) => 
                           AND_OUT_17_port, OUT_LOGIC_AND(16) => 
                           AND_OUT_16_port, OUT_LOGIC_AND(15) => 
                           AND_OUT_15_port, OUT_LOGIC_AND(14) => 
                           AND_OUT_14_port, OUT_LOGIC_AND(13) => 
                           AND_OUT_13_port, OUT_LOGIC_AND(12) => 
                           AND_OUT_12_port, OUT_LOGIC_AND(11) => 
                           AND_OUT_11_port, OUT_LOGIC_AND(10) => 
                           AND_OUT_10_port, OUT_LOGIC_AND(9) => AND_OUT_9_port,
                           OUT_LOGIC_AND(8) => AND_OUT_8_port, OUT_LOGIC_AND(7)
                           => AND_OUT_7_port, OUT_LOGIC_AND(6) => 
                           AND_OUT_6_port, OUT_LOGIC_AND(5) => AND_OUT_5_port, 
                           OUT_LOGIC_AND(4) => AND_OUT_4_port, OUT_LOGIC_AND(3)
                           => AND_OUT_3_port, OUT_LOGIC_AND(2) => 
                           AND_OUT_2_port, OUT_LOGIC_AND(1) => AND_OUT_1_port, 
                           OUT_LOGIC_AND(0) => AND_OUT_0_port, OUT_LOGIC_OR(31)
                           => OR_OUT_31_port, OUT_LOGIC_OR(30) => 
                           OR_OUT_30_port, OUT_LOGIC_OR(29) => OR_OUT_29_port, 
                           OUT_LOGIC_OR(28) => OR_OUT_28_port, OUT_LOGIC_OR(27)
                           => OR_OUT_27_port, OUT_LOGIC_OR(26) => 
                           OR_OUT_26_port, OUT_LOGIC_OR(25) => OR_OUT_25_port, 
                           OUT_LOGIC_OR(24) => OR_OUT_24_port, OUT_LOGIC_OR(23)
                           => OR_OUT_23_port, OUT_LOGIC_OR(22) => 
                           OR_OUT_22_port, OUT_LOGIC_OR(21) => OR_OUT_21_port, 
                           OUT_LOGIC_OR(20) => OR_OUT_20_port, OUT_LOGIC_OR(19)
                           => OR_OUT_19_port, OUT_LOGIC_OR(18) => 
                           OR_OUT_18_port, OUT_LOGIC_OR(17) => OR_OUT_17_port, 
                           OUT_LOGIC_OR(16) => OR_OUT_16_port, OUT_LOGIC_OR(15)
                           => OR_OUT_15_port, OUT_LOGIC_OR(14) => 
                           OR_OUT_14_port, OUT_LOGIC_OR(13) => OR_OUT_13_port, 
                           OUT_LOGIC_OR(12) => OR_OUT_12_port, OUT_LOGIC_OR(11)
                           => OR_OUT_11_port, OUT_LOGIC_OR(10) => 
                           OR_OUT_10_port, OUT_LOGIC_OR(9) => OR_OUT_9_port, 
                           OUT_LOGIC_OR(8) => OR_OUT_8_port, OUT_LOGIC_OR(7) =>
                           OR_OUT_7_port, OUT_LOGIC_OR(6) => OR_OUT_6_port, 
                           OUT_LOGIC_OR(5) => OR_OUT_5_port, OUT_LOGIC_OR(4) =>
                           OR_OUT_4_port, OUT_LOGIC_OR(3) => OR_OUT_3_port, 
                           OUT_LOGIC_OR(2) => OR_OUT_2_port, OUT_LOGIC_OR(1) =>
                           OR_OUT_1_port, OUT_LOGIC_OR(0) => OR_OUT_0_port, 
                           OUT_LOGIC_XOR(31) => XOR_OUT_31_port, 
                           OUT_LOGIC_XOR(30) => XOR_OUT_30_port, 
                           OUT_LOGIC_XOR(29) => XOR_OUT_29_port, 
                           OUT_LOGIC_XOR(28) => XOR_OUT_28_port, 
                           OUT_LOGIC_XOR(27) => XOR_OUT_27_port, 
                           OUT_LOGIC_XOR(26) => XOR_OUT_26_port, 
                           OUT_LOGIC_XOR(25) => XOR_OUT_25_port, 
                           OUT_LOGIC_XOR(24) => XOR_OUT_24_port, 
                           OUT_LOGIC_XOR(23) => XOR_OUT_23_port, 
                           OUT_LOGIC_XOR(22) => XOR_OUT_22_port, 
                           OUT_LOGIC_XOR(21) => XOR_OUT_21_port, 
                           OUT_LOGIC_XOR(20) => XOR_OUT_20_port, 
                           OUT_LOGIC_XOR(19) => XOR_OUT_19_port, 
                           OUT_LOGIC_XOR(18) => XOR_OUT_18_port, 
                           OUT_LOGIC_XOR(17) => XOR_OUT_17_port, 
                           OUT_LOGIC_XOR(16) => XOR_OUT_16_port, 
                           OUT_LOGIC_XOR(15) => XOR_OUT_15_port, 
                           OUT_LOGIC_XOR(14) => XOR_OUT_14_port, 
                           OUT_LOGIC_XOR(13) => XOR_OUT_13_port, 
                           OUT_LOGIC_XOR(12) => XOR_OUT_12_port, 
                           OUT_LOGIC_XOR(11) => XOR_OUT_11_port, 
                           OUT_LOGIC_XOR(10) => XOR_OUT_10_port, 
                           OUT_LOGIC_XOR(9) => XOR_OUT_9_port, OUT_LOGIC_XOR(8)
                           => XOR_OUT_8_port, OUT_LOGIC_XOR(7) => 
                           XOR_OUT_7_port, OUT_LOGIC_XOR(6) => XOR_OUT_6_port, 
                           OUT_LOGIC_XOR(5) => XOR_OUT_5_port, OUT_LOGIC_XOR(4)
                           => XOR_OUT_4_port, OUT_LOGIC_XOR(3) => 
                           XOR_OUT_3_port, OUT_LOGIC_XOR(2) => XOR_OUT_2_port, 
                           OUT_LOGIC_XOR(1) => XOR_OUT_1_port, OUT_LOGIC_XOR(0)
                           => XOR_OUT_0_port);
   adder_sub : p4_adder_N32_N_carry4 port map( A(31) => DATA1(31), A(30) => 
                           DATA1(30), A(29) => DATA1(29), A(28) => DATA1(28), 
                           A(27) => DATA1(27), A(26) => DATA1(26), A(25) => 
                           DATA1(25), A(24) => DATA1(24), A(23) => DATA1(23), 
                           A(22) => DATA1(22), A(21) => DATA1(21), A(20) => 
                           DATA1(20), A(19) => DATA1(19), A(18) => DATA1(18), 
                           A(17) => DATA1(17), A(16) => DATA1(16), A(15) => 
                           DATA1(15), A(14) => DATA1(14), A(13) => DATA1(13), 
                           A(12) => DATA1(12), A(11) => DATA1(11), A(10) => 
                           DATA1(10), A(9) => DATA1(9), A(8) => DATA1(8), A(7) 
                           => DATA1(7), A(6) => DATA1(6), A(5) => DATA1(5), 
                           A(4) => DATA1(4), A(3) => DATA1(3), A(2) => DATA1(2)
                           , A(1) => DATA1(1), A(0) => DATA1(0), B(31) => 
                           DATA2(31), B(30) => DATA2(30), B(29) => DATA2(29), 
                           B(28) => DATA2(28), B(27) => DATA2(27), B(26) => 
                           DATA2(26), B(25) => DATA2(25), B(24) => DATA2(24), 
                           B(23) => DATA2(23), B(22) => DATA2(22), B(21) => 
                           DATA2(21), B(20) => DATA2(20), B(19) => DATA2(19), 
                           B(18) => DATA2(18), B(17) => DATA2(17), B(16) => 
                           DATA2(16), B(15) => DATA2(15), B(14) => DATA2(14), 
                           B(13) => DATA2(13), B(12) => DATA2(12), B(11) => 
                           DATA2(11), B(10) => DATA2(10), B(9) => DATA2(9), 
                           B(8) => DATA2(8), B(7) => DATA2(7), B(6) => DATA2(6)
                           , B(5) => DATA2(5), B(4) => DATA2(4), B(3) => 
                           DATA2(3), B(2) => DATA2(2), B(1) => DATA2(1), B(0) 
                           => DATA2(0), Cin => Add_subn, SUM(31) => 
                           add_sub_out_31_port, SUM(30) => add_sub_out_30_port,
                           SUM(29) => add_sub_out_29_port, SUM(28) => 
                           add_sub_out_28_port, SUM(27) => add_sub_out_27_port,
                           SUM(26) => add_sub_out_26_port, SUM(25) => 
                           add_sub_out_25_port, SUM(24) => add_sub_out_24_port,
                           SUM(23) => add_sub_out_23_port, SUM(22) => 
                           add_sub_out_22_port, SUM(21) => add_sub_out_21_port,
                           SUM(20) => add_sub_out_20_port, SUM(19) => 
                           add_sub_out_19_port, SUM(18) => add_sub_out_18_port,
                           SUM(17) => add_sub_out_17_port, SUM(16) => 
                           add_sub_out_16_port, SUM(15) => add_sub_out_15_port,
                           SUM(14) => add_sub_out_14_port, SUM(13) => 
                           add_sub_out_13_port, SUM(12) => add_sub_out_12_port,
                           SUM(11) => add_sub_out_11_port, SUM(10) => 
                           add_sub_out_10_port, SUM(9) => add_sub_out_9_port, 
                           SUM(8) => add_sub_out_8_port, SUM(7) => 
                           add_sub_out_7_port, SUM(6) => add_sub_out_6_port, 
                           SUM(5) => add_sub_out_5_port, SUM(4) => 
                           add_sub_out_4_port, SUM(3) => add_sub_out_3_port, 
                           SUM(2) => add_sub_out_2_port, SUM(1) => 
                           add_sub_out_1_port, SUM(0) => add_sub_out_0_port);
   comp : compare_N32 port map( num1(31) => DATA1(31), num1(30) => DATA1(30), 
                           num1(29) => DATA1(29), num1(28) => DATA1(28), 
                           num1(27) => DATA1(27), num1(26) => DATA1(26), 
                           num1(25) => DATA1(25), num1(24) => DATA1(24), 
                           num1(23) => DATA1(23), num1(22) => DATA1(22), 
                           num1(21) => DATA1(21), num1(20) => DATA1(20), 
                           num1(19) => DATA1(19), num1(18) => DATA1(18), 
                           num1(17) => DATA1(17), num1(16) => DATA1(16), 
                           num1(15) => DATA1(15), num1(14) => DATA1(14), 
                           num1(13) => DATA1(13), num1(12) => DATA1(12), 
                           num1(11) => DATA1(11), num1(10) => DATA1(10), 
                           num1(9) => DATA1(9), num1(8) => DATA1(8), num1(7) =>
                           DATA1(7), num1(6) => DATA1(6), num1(5) => DATA1(5), 
                           num1(4) => DATA1(4), num1(3) => DATA1(3), num1(2) =>
                           DATA1(2), num1(1) => DATA1(1), num1(0) => DATA1(0), 
                           num2(31) => DATA2(31), num2(30) => DATA2(30), 
                           num2(29) => DATA2(29), num2(28) => DATA2(28), 
                           num2(27) => DATA2(27), num2(26) => DATA2(26), 
                           num2(25) => DATA2(25), num2(24) => DATA2(24), 
                           num2(23) => DATA2(23), num2(22) => DATA2(22), 
                           num2(21) => DATA2(21), num2(20) => DATA2(20), 
                           num2(19) => DATA2(19), num2(18) => DATA2(18), 
                           num2(17) => DATA2(17), num2(16) => DATA2(16), 
                           num2(15) => DATA2(15), num2(14) => DATA2(14), 
                           num2(13) => DATA2(13), num2(12) => DATA2(12), 
                           num2(11) => DATA2(11), num2(10) => DATA2(10), 
                           num2(9) => DATA2(9), num2(8) => DATA2(8), num2(7) =>
                           DATA2(7), num2(6) => DATA2(6), num2(5) => DATA2(5), 
                           num2(4) => DATA2(4), num2(3) => DATA2(3), num2(2) =>
                           DATA2(2), num2(1) => DATA2(1), num2(0) => DATA2(0), 
                           less => net2103, equal => comp_eq, greater => 
                           comp_greater);
   mux_comp : MUX_2to1_n32 port map( A(31) => X_Logic0_port, A(30) => 
                           X_Logic0_port, A(29) => X_Logic0_port, A(28) => 
                           X_Logic0_port, A(27) => X_Logic0_port, A(26) => 
                           X_Logic0_port, A(25) => X_Logic0_port, A(24) => 
                           X_Logic0_port, A(23) => X_Logic0_port, A(22) => 
                           X_Logic0_port, A(21) => X_Logic0_port, A(20) => 
                           X_Logic0_port, A(19) => X_Logic0_port, A(18) => 
                           X_Logic0_port, A(17) => X_Logic0_port, A(16) => 
                           X_Logic0_port, A(15) => X_Logic0_port, A(14) => 
                           X_Logic0_port, A(13) => X_Logic0_port, A(12) => 
                           X_Logic0_port, A(11) => X_Logic0_port, A(10) => 
                           X_Logic0_port, A(9) => X_Logic0_port, A(8) => 
                           X_Logic0_port, A(7) => X_Logic0_port, A(6) => 
                           X_Logic0_port, A(5) => X_Logic0_port, A(4) => 
                           X_Logic0_port, A(3) => X_Logic0_port, A(2) => 
                           X_Logic0_port, A(1) => X_Logic0_port, A(0) => 
                           X_Logic0_port, B(31) => X_Logic0_port, B(30) => 
                           X_Logic0_port, B(29) => X_Logic0_port, B(28) => 
                           X_Logic0_port, B(27) => X_Logic0_port, B(26) => 
                           X_Logic0_port, B(25) => X_Logic0_port, B(24) => 
                           X_Logic0_port, B(23) => X_Logic0_port, B(22) => 
                           X_Logic0_port, B(21) => X_Logic0_port, B(20) => 
                           X_Logic0_port, B(19) => X_Logic0_port, B(18) => 
                           X_Logic0_port, B(17) => X_Logic0_port, B(16) => 
                           X_Logic0_port, B(15) => X_Logic0_port, B(14) => 
                           X_Logic0_port, B(13) => X_Logic0_port, B(12) => 
                           X_Logic0_port, B(11) => X_Logic0_port, B(10) => 
                           X_Logic0_port, B(9) => X_Logic0_port, B(8) => 
                           X_Logic0_port, B(7) => X_Logic0_port, B(6) => 
                           X_Logic0_port, B(5) => X_Logic0_port, B(4) => 
                           X_Logic0_port, B(3) => X_Logic0_port, B(2) => 
                           X_Logic0_port, B(1) => X_Logic0_port, B(0) => 
                           X_Logic1_port, S => sel_mux_comp_out, Y(31) => 
                           comp_out_31_port, Y(30) => comp_out_30_port, Y(29) 
                           => comp_out_29_port, Y(28) => comp_out_28_port, 
                           Y(27) => comp_out_27_port, Y(26) => comp_out_26_port
                           , Y(25) => comp_out_25_port, Y(24) => 
                           comp_out_24_port, Y(23) => comp_out_23_port, Y(22) 
                           => comp_out_22_port, Y(21) => comp_out_21_port, 
                           Y(20) => comp_out_20_port, Y(19) => comp_out_19_port
                           , Y(18) => comp_out_18_port, Y(17) => 
                           comp_out_17_port, Y(16) => comp_out_16_port, Y(15) 
                           => comp_out_15_port, Y(14) => comp_out_14_port, 
                           Y(13) => comp_out_13_port, Y(12) => comp_out_12_port
                           , Y(11) => comp_out_11_port, Y(10) => 
                           comp_out_10_port, Y(9) => comp_out_9_port, Y(8) => 
                           comp_out_8_port, Y(7) => comp_out_7_port, Y(6) => 
                           comp_out_6_port, Y(5) => comp_out_5_port, Y(4) => 
                           comp_out_4_port, Y(3) => comp_out_3_port, Y(2) => 
                           comp_out_2_port, Y(1) => comp_out_1_port, Y(0) => 
                           comp_out_0_port);
   mux_alu_out : MUX_6to1_n32 port map( A(31) => add_sub_out_31_port, A(30) => 
                           add_sub_out_30_port, A(29) => add_sub_out_29_port, 
                           A(28) => add_sub_out_28_port, A(27) => 
                           add_sub_out_27_port, A(26) => add_sub_out_26_port, 
                           A(25) => add_sub_out_25_port, A(24) => 
                           add_sub_out_24_port, A(23) => add_sub_out_23_port, 
                           A(22) => add_sub_out_22_port, A(21) => 
                           add_sub_out_21_port, A(20) => add_sub_out_20_port, 
                           A(19) => add_sub_out_19_port, A(18) => 
                           add_sub_out_18_port, A(17) => add_sub_out_17_port, 
                           A(16) => add_sub_out_16_port, A(15) => 
                           add_sub_out_15_port, A(14) => add_sub_out_14_port, 
                           A(13) => add_sub_out_13_port, A(12) => 
                           add_sub_out_12_port, A(11) => add_sub_out_11_port, 
                           A(10) => add_sub_out_10_port, A(9) => 
                           add_sub_out_9_port, A(8) => add_sub_out_8_port, A(7)
                           => add_sub_out_7_port, A(6) => add_sub_out_6_port, 
                           A(5) => add_sub_out_5_port, A(4) => 
                           add_sub_out_4_port, A(3) => add_sub_out_3_port, A(2)
                           => add_sub_out_2_port, A(1) => add_sub_out_1_port, 
                           A(0) => add_sub_out_0_port, B(31) => AND_OUT_31_port
                           , B(30) => AND_OUT_30_port, B(29) => AND_OUT_29_port
                           , B(28) => AND_OUT_28_port, B(27) => AND_OUT_27_port
                           , B(26) => AND_OUT_26_port, B(25) => AND_OUT_25_port
                           , B(24) => AND_OUT_24_port, B(23) => AND_OUT_23_port
                           , B(22) => AND_OUT_22_port, B(21) => AND_OUT_21_port
                           , B(20) => AND_OUT_20_port, B(19) => AND_OUT_19_port
                           , B(18) => AND_OUT_18_port, B(17) => AND_OUT_17_port
                           , B(16) => AND_OUT_16_port, B(15) => AND_OUT_15_port
                           , B(14) => AND_OUT_14_port, B(13) => AND_OUT_13_port
                           , B(12) => AND_OUT_12_port, B(11) => AND_OUT_11_port
                           , B(10) => AND_OUT_10_port, B(9) => AND_OUT_9_port, 
                           B(8) => AND_OUT_8_port, B(7) => AND_OUT_7_port, B(6)
                           => AND_OUT_6_port, B(5) => AND_OUT_5_port, B(4) => 
                           AND_OUT_4_port, B(3) => AND_OUT_3_port, B(2) => 
                           AND_OUT_2_port, B(1) => AND_OUT_1_port, B(0) => 
                           AND_OUT_0_port, C(31) => OR_OUT_31_port, C(30) => 
                           OR_OUT_30_port, C(29) => OR_OUT_29_port, C(28) => 
                           OR_OUT_28_port, C(27) => OR_OUT_27_port, C(26) => 
                           OR_OUT_26_port, C(25) => OR_OUT_25_port, C(24) => 
                           OR_OUT_24_port, C(23) => OR_OUT_23_port, C(22) => 
                           OR_OUT_22_port, C(21) => OR_OUT_21_port, C(20) => 
                           OR_OUT_20_port, C(19) => OR_OUT_19_port, C(18) => 
                           OR_OUT_18_port, C(17) => OR_OUT_17_port, C(16) => 
                           OR_OUT_16_port, C(15) => OR_OUT_15_port, C(14) => 
                           OR_OUT_14_port, C(13) => OR_OUT_13_port, C(12) => 
                           OR_OUT_12_port, C(11) => OR_OUT_11_port, C(10) => 
                           OR_OUT_10_port, C(9) => OR_OUT_9_port, C(8) => 
                           OR_OUT_8_port, C(7) => OR_OUT_7_port, C(6) => 
                           OR_OUT_6_port, C(5) => OR_OUT_5_port, C(4) => 
                           OR_OUT_4_port, C(3) => OR_OUT_3_port, C(2) => 
                           OR_OUT_2_port, C(1) => OR_OUT_1_port, C(0) => 
                           OR_OUT_0_port, D(31) => XOR_OUT_31_port, D(30) => 
                           XOR_OUT_30_port, D(29) => XOR_OUT_29_port, D(28) => 
                           XOR_OUT_28_port, D(27) => XOR_OUT_27_port, D(26) => 
                           XOR_OUT_26_port, D(25) => XOR_OUT_25_port, D(24) => 
                           XOR_OUT_24_port, D(23) => XOR_OUT_23_port, D(22) => 
                           XOR_OUT_22_port, D(21) => XOR_OUT_21_port, D(20) => 
                           XOR_OUT_20_port, D(19) => XOR_OUT_19_port, D(18) => 
                           XOR_OUT_18_port, D(17) => XOR_OUT_17_port, D(16) => 
                           XOR_OUT_16_port, D(15) => XOR_OUT_15_port, D(14) => 
                           XOR_OUT_14_port, D(13) => XOR_OUT_13_port, D(12) => 
                           XOR_OUT_12_port, D(11) => XOR_OUT_11_port, D(10) => 
                           XOR_OUT_10_port, D(9) => XOR_OUT_9_port, D(8) => 
                           XOR_OUT_8_port, D(7) => XOR_OUT_7_port, D(6) => 
                           XOR_OUT_6_port, D(5) => XOR_OUT_5_port, D(4) => 
                           XOR_OUT_4_port, D(3) => XOR_OUT_3_port, D(2) => 
                           XOR_OUT_2_port, D(1) => XOR_OUT_1_port, D(0) => 
                           XOR_OUT_0_port, E(31) => comp_out_31_port, E(30) => 
                           comp_out_30_port, E(29) => comp_out_29_port, E(28) 
                           => comp_out_28_port, E(27) => comp_out_27_port, 
                           E(26) => comp_out_26_port, E(25) => comp_out_25_port
                           , E(24) => comp_out_24_port, E(23) => 
                           comp_out_23_port, E(22) => comp_out_22_port, E(21) 
                           => comp_out_21_port, E(20) => comp_out_20_port, 
                           E(19) => comp_out_19_port, E(18) => comp_out_18_port
                           , E(17) => comp_out_17_port, E(16) => 
                           comp_out_16_port, E(15) => comp_out_15_port, E(14) 
                           => comp_out_14_port, E(13) => comp_out_13_port, 
                           E(12) => comp_out_12_port, E(11) => comp_out_11_port
                           , E(10) => comp_out_10_port, E(9) => comp_out_9_port
                           , E(8) => comp_out_8_port, E(7) => comp_out_7_port, 
                           E(6) => comp_out_6_port, E(5) => comp_out_5_port, 
                           E(4) => comp_out_4_port, E(3) => comp_out_3_port, 
                           E(2) => comp_out_2_port, E(1) => comp_out_1_port, 
                           E(0) => comp_out_0_port, F(31) => shift_out_31_port,
                           F(30) => shift_out_30_port, F(29) => 
                           shift_out_29_port, F(28) => shift_out_28_port, F(27)
                           => shift_out_27_port, F(26) => shift_out_26_port, 
                           F(25) => shift_out_25_port, F(24) => 
                           shift_out_24_port, F(23) => shift_out_23_port, F(22)
                           => shift_out_22_port, F(21) => shift_out_21_port, 
                           F(20) => shift_out_20_port, F(19) => 
                           shift_out_19_port, F(18) => shift_out_18_port, F(17)
                           => shift_out_17_port, F(16) => shift_out_16_port, 
                           F(15) => shift_out_15_port, F(14) => 
                           shift_out_14_port, F(13) => shift_out_13_port, F(12)
                           => shift_out_12_port, F(11) => shift_out_11_port, 
                           F(10) => shift_out_10_port, F(9) => shift_out_9_port
                           , F(8) => shift_out_8_port, F(7) => shift_out_7_port
                           , F(6) => shift_out_6_port, F(5) => shift_out_5_port
                           , F(4) => shift_out_4_port, F(3) => shift_out_3_port
                           , F(2) => shift_out_2_port, F(1) => shift_out_1_port
                           , F(0) => shift_out_0_port, S(2) => AluOpCode(2), 
                           S(1) => AluOpCode(1), S(0) => AluOpCode(0), Y(31) =>
                           OUTALU(31), Y(30) => OUTALU(30), Y(29) => OUTALU(29)
                           , Y(28) => OUTALU(28), Y(27) => OUTALU(27), Y(26) =>
                           OUTALU(26), Y(25) => OUTALU(25), Y(24) => OUTALU(24)
                           , Y(23) => OUTALU(23), Y(22) => OUTALU(22), Y(21) =>
                           OUTALU(21), Y(20) => OUTALU(20), Y(19) => OUTALU(19)
                           , Y(18) => OUTALU(18), Y(17) => OUTALU(17), Y(16) =>
                           OUTALU(16), Y(15) => OUTALU(15), Y(14) => OUTALU(14)
                           , Y(13) => OUTALU(13), Y(12) => OUTALU(12), Y(11) =>
                           OUTALU(11), Y(10) => OUTALU(10), Y(9) => OUTALU(9), 
                           Y(8) => OUTALU(8), Y(7) => OUTALU(7), Y(6) => 
                           OUTALU(6), Y(5) => OUTALU(5), Y(4) => OUTALU(4), 
                           Y(3) => OUTALU(3), Y(2) => OUTALU(2), Y(1) => 
                           OUTALU(1), Y(0) => OUTALU(0));
   U3 : NAND2_X2 port map( A1 => n1, A2 => n2, ZN => sel_mux_comp_out);
   U4 : OAI21_X1 port map( B1 => comp_eq, B2 => comp_greater, A => 
                           CompareOpCode(1), ZN => n2);
   U5 : NAND2_X1 port map( A1 => CompareOpCode(0), A2 => n3, ZN => n1);
   U6 : INV_X1 port map( A => comp_eq, ZN => n3);
   U7 : MUX2_X1 port map( A => CompareOpCode(2), B => CompareOpCode(3), S => 
                           comp_eq, Z => CompBranch);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N5_0 is

   port( data : in std_logic_vector (4 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (4 downto 0));

end registro_N5_0;

architecture SYN_behaviour of registro_N5_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n11, n12, n13, n14,
      n15, net43246, net43247, net43248, net43249, net43250 : std_logic;

begin
   Q <= ( Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_4_inst : DFFR_X1 port map( D => n15, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43250);
   Q_reg_3_inst : DFFR_X1 port map( D => n14, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43249);
   Q_reg_2_inst : DFFR_X1 port map( D => n13, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43248);
   Q_reg_1_inst : DFFR_X1 port map( D => n12, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43247);
   Q_reg_0_inst : DFFR_X1 port map( D => n11, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43246);
   U2 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n15);
   U3 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n14);
   U4 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n13);
   U5 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n12);
   U6 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n11);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N17 is

   port( data : in std_logic_vector (16 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (16 downto 0));

end registro_N17;

architecture SYN_behaviour of registro_N17 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_16_port, Q_15_port, Q_14_port, Q_13_port, Q_12_port, Q_11_port, 
      Q_10_port, Q_9_port, Q_8_port, Q_7_port, Q_6_port, Q_5_port, Q_4_port, 
      Q_3_port, Q_2_port, Q_1_port, Q_0_port, n35, n36, n37, n38, n39, n40, n41
      , n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, net43229, net43230, 
      net43231, net43232, net43233, net43234, net43235, net43236, net43237, 
      net43238, net43239, net43240, net43241, net43242, net43243, net43244, 
      net43245 : std_logic;

begin
   Q <= ( Q_16_port, Q_15_port, Q_14_port, Q_13_port, Q_12_port, Q_11_port, 
      Q_10_port, Q_9_port, Q_8_port, Q_7_port, Q_6_port, Q_5_port, Q_4_port, 
      Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_16_inst : DFFR_X1 port map( D => n51, CK => clock, RN => clear, Q => 
                           Q_16_port, QN => net43245);
   Q_reg_15_inst : DFFR_X1 port map( D => n50, CK => clock, RN => clear, Q => 
                           Q_15_port, QN => net43244);
   Q_reg_14_inst : DFFR_X1 port map( D => n49, CK => clock, RN => clear, Q => 
                           Q_14_port, QN => net43243);
   Q_reg_13_inst : DFFR_X1 port map( D => n48, CK => clock, RN => clear, Q => 
                           Q_13_port, QN => net43242);
   Q_reg_12_inst : DFFR_X1 port map( D => n47, CK => clock, RN => clear, Q => 
                           Q_12_port, QN => net43241);
   Q_reg_11_inst : DFFR_X1 port map( D => n46, CK => clock, RN => clear, Q => 
                           Q_11_port, QN => net43240);
   Q_reg_10_inst : DFFR_X1 port map( D => n45, CK => clock, RN => clear, Q => 
                           Q_10_port, QN => net43239);
   Q_reg_9_inst : DFFR_X1 port map( D => n44, CK => clock, RN => clear, Q => 
                           Q_9_port, QN => net43238);
   Q_reg_8_inst : DFFR_X1 port map( D => n43, CK => clock, RN => clear, Q => 
                           Q_8_port, QN => net43237);
   Q_reg_7_inst : DFFR_X1 port map( D => n42, CK => clock, RN => clear, Q => 
                           Q_7_port, QN => net43236);
   Q_reg_6_inst : DFFR_X1 port map( D => n41, CK => clock, RN => clear, Q => 
                           Q_6_port, QN => net43235);
   Q_reg_5_inst : DFFR_X1 port map( D => n40, CK => clock, RN => clear, Q => 
                           Q_5_port, QN => net43234);
   Q_reg_4_inst : DFFR_X1 port map( D => n39, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43233);
   Q_reg_3_inst : DFFR_X1 port map( D => n38, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43232);
   Q_reg_2_inst : DFFR_X1 port map( D => n37, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43231);
   Q_reg_1_inst : DFFR_X1 port map( D => n36, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43230);
   Q_reg_0_inst : DFFR_X1 port map( D => n35, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43229);
   U2 : MUX2_X1 port map( A => Q_16_port, B => data(16), S => enable, Z => n51)
                           ;
   U3 : MUX2_X1 port map( A => Q_15_port, B => data(15), S => enable, Z => n50)
                           ;
   U4 : MUX2_X1 port map( A => Q_14_port, B => data(14), S => enable, Z => n49)
                           ;
   U5 : MUX2_X1 port map( A => Q_13_port, B => data(13), S => enable, Z => n48)
                           ;
   U6 : MUX2_X1 port map( A => Q_12_port, B => data(12), S => enable, Z => n47)
                           ;
   U7 : MUX2_X1 port map( A => Q_11_port, B => data(11), S => enable, Z => n46)
                           ;
   U8 : MUX2_X1 port map( A => Q_10_port, B => data(10), S => enable, Z => n45)
                           ;
   U9 : MUX2_X1 port map( A => Q_9_port, B => data(9), S => enable, Z => n44);
   U10 : MUX2_X1 port map( A => Q_8_port, B => data(8), S => enable, Z => n43);
   U11 : MUX2_X1 port map( A => Q_7_port, B => data(7), S => enable, Z => n42);
   U12 : MUX2_X1 port map( A => Q_6_port, B => data(6), S => enable, Z => n41);
   U13 : MUX2_X1 port map( A => Q_5_port, B => data(5), S => enable, Z => n40);
   U14 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n39);
   U15 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n38);
   U16 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n37);
   U17 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n36);
   U18 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n35);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity registro_N32_0 is

   port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : in 
         std_logic;  Q : out std_logic_vector (31 downto 0));

end registro_N32_0;

architecture SYN_behaviour of registro_N32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port, n65
      , n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, 
      n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94
      , n95, n96, net43197, net43198, net43199, net43200, net43201, net43202, 
      net43203, net43204, net43205, net43206, net43207, net43208, net43209, 
      net43210, net43211, net43212, net43213, net43214, net43215, net43216, 
      net43217, net43218, net43219, net43220, net43221, net43222, net43223, 
      net43224, net43225, net43226, net43227, net43228 : std_logic;

begin
   Q <= ( Q_31_port, Q_30_port, Q_29_port, Q_28_port, Q_27_port, Q_26_port, 
      Q_25_port, Q_24_port, Q_23_port, Q_22_port, Q_21_port, Q_20_port, 
      Q_19_port, Q_18_port, Q_17_port, Q_16_port, Q_15_port, Q_14_port, 
      Q_13_port, Q_12_port, Q_11_port, Q_10_port, Q_9_port, Q_8_port, Q_7_port,
      Q_6_port, Q_5_port, Q_4_port, Q_3_port, Q_2_port, Q_1_port, Q_0_port );
   
   Q_reg_31_inst : DFFR_X1 port map( D => n96, CK => clock, RN => clear, Q => 
                           Q_31_port, QN => net43228);
   Q_reg_30_inst : DFFR_X1 port map( D => n95, CK => clock, RN => clear, Q => 
                           Q_30_port, QN => net43227);
   Q_reg_29_inst : DFFR_X1 port map( D => n94, CK => clock, RN => clear, Q => 
                           Q_29_port, QN => net43226);
   Q_reg_28_inst : DFFR_X1 port map( D => n93, CK => clock, RN => clear, Q => 
                           Q_28_port, QN => net43225);
   Q_reg_27_inst : DFFR_X1 port map( D => n92, CK => clock, RN => clear, Q => 
                           Q_27_port, QN => net43224);
   Q_reg_26_inst : DFFR_X1 port map( D => n91, CK => clock, RN => clear, Q => 
                           Q_26_port, QN => net43223);
   Q_reg_25_inst : DFFR_X1 port map( D => n90, CK => clock, RN => clear, Q => 
                           Q_25_port, QN => net43222);
   Q_reg_24_inst : DFFR_X1 port map( D => n89, CK => clock, RN => clear, Q => 
                           Q_24_port, QN => net43221);
   Q_reg_23_inst : DFFR_X1 port map( D => n88, CK => clock, RN => clear, Q => 
                           Q_23_port, QN => net43220);
   Q_reg_22_inst : DFFR_X1 port map( D => n87, CK => clock, RN => clear, Q => 
                           Q_22_port, QN => net43219);
   Q_reg_21_inst : DFFR_X1 port map( D => n86, CK => clock, RN => clear, Q => 
                           Q_21_port, QN => net43218);
   Q_reg_20_inst : DFFR_X1 port map( D => n85, CK => clock, RN => clear, Q => 
                           Q_20_port, QN => net43217);
   Q_reg_19_inst : DFFR_X1 port map( D => n84, CK => clock, RN => clear, Q => 
                           Q_19_port, QN => net43216);
   Q_reg_18_inst : DFFR_X1 port map( D => n83, CK => clock, RN => clear, Q => 
                           Q_18_port, QN => net43215);
   Q_reg_17_inst : DFFR_X1 port map( D => n82, CK => clock, RN => clear, Q => 
                           Q_17_port, QN => net43214);
   Q_reg_16_inst : DFFR_X1 port map( D => n81, CK => clock, RN => clear, Q => 
                           Q_16_port, QN => net43213);
   Q_reg_15_inst : DFFR_X1 port map( D => n80, CK => clock, RN => clear, Q => 
                           Q_15_port, QN => net43212);
   Q_reg_14_inst : DFFR_X1 port map( D => n79, CK => clock, RN => clear, Q => 
                           Q_14_port, QN => net43211);
   Q_reg_13_inst : DFFR_X1 port map( D => n78, CK => clock, RN => clear, Q => 
                           Q_13_port, QN => net43210);
   Q_reg_12_inst : DFFR_X1 port map( D => n77, CK => clock, RN => clear, Q => 
                           Q_12_port, QN => net43209);
   Q_reg_11_inst : DFFR_X1 port map( D => n76, CK => clock, RN => clear, Q => 
                           Q_11_port, QN => net43208);
   Q_reg_10_inst : DFFR_X1 port map( D => n75, CK => clock, RN => clear, Q => 
                           Q_10_port, QN => net43207);
   Q_reg_9_inst : DFFR_X1 port map( D => n74, CK => clock, RN => clear, Q => 
                           Q_9_port, QN => net43206);
   Q_reg_8_inst : DFFR_X1 port map( D => n73, CK => clock, RN => clear, Q => 
                           Q_8_port, QN => net43205);
   Q_reg_7_inst : DFFR_X1 port map( D => n72, CK => clock, RN => clear, Q => 
                           Q_7_port, QN => net43204);
   Q_reg_6_inst : DFFR_X1 port map( D => n71, CK => clock, RN => clear, Q => 
                           Q_6_port, QN => net43203);
   Q_reg_5_inst : DFFR_X1 port map( D => n70, CK => clock, RN => clear, Q => 
                           Q_5_port, QN => net43202);
   Q_reg_4_inst : DFFR_X1 port map( D => n69, CK => clock, RN => clear, Q => 
                           Q_4_port, QN => net43201);
   Q_reg_3_inst : DFFR_X1 port map( D => n68, CK => clock, RN => clear, Q => 
                           Q_3_port, QN => net43200);
   Q_reg_2_inst : DFFR_X1 port map( D => n67, CK => clock, RN => clear, Q => 
                           Q_2_port, QN => net43199);
   Q_reg_1_inst : DFFR_X1 port map( D => n66, CK => clock, RN => clear, Q => 
                           Q_1_port, QN => net43198);
   Q_reg_0_inst : DFFR_X1 port map( D => n65, CK => clock, RN => clear, Q => 
                           Q_0_port, QN => net43197);
   U2 : MUX2_X1 port map( A => Q_31_port, B => data(31), S => enable, Z => n96)
                           ;
   U3 : MUX2_X1 port map( A => Q_30_port, B => data(30), S => enable, Z => n95)
                           ;
   U4 : MUX2_X1 port map( A => Q_29_port, B => data(29), S => enable, Z => n94)
                           ;
   U5 : MUX2_X1 port map( A => Q_28_port, B => data(28), S => enable, Z => n93)
                           ;
   U6 : MUX2_X1 port map( A => Q_27_port, B => data(27), S => enable, Z => n92)
                           ;
   U7 : MUX2_X1 port map( A => Q_26_port, B => data(26), S => enable, Z => n91)
                           ;
   U8 : MUX2_X1 port map( A => Q_25_port, B => data(25), S => enable, Z => n90)
                           ;
   U9 : MUX2_X1 port map( A => Q_24_port, B => data(24), S => enable, Z => n89)
                           ;
   U10 : MUX2_X1 port map( A => Q_23_port, B => data(23), S => enable, Z => n88
                           );
   U11 : MUX2_X1 port map( A => Q_22_port, B => data(22), S => enable, Z => n87
                           );
   U12 : MUX2_X1 port map( A => Q_21_port, B => data(21), S => enable, Z => n86
                           );
   U13 : MUX2_X1 port map( A => Q_20_port, B => data(20), S => enable, Z => n85
                           );
   U14 : MUX2_X1 port map( A => Q_19_port, B => data(19), S => enable, Z => n84
                           );
   U15 : MUX2_X1 port map( A => Q_18_port, B => data(18), S => enable, Z => n83
                           );
   U16 : MUX2_X1 port map( A => Q_17_port, B => data(17), S => enable, Z => n82
                           );
   U17 : MUX2_X1 port map( A => Q_16_port, B => data(16), S => enable, Z => n81
                           );
   U18 : MUX2_X1 port map( A => Q_15_port, B => data(15), S => enable, Z => n80
                           );
   U19 : MUX2_X1 port map( A => Q_14_port, B => data(14), S => enable, Z => n79
                           );
   U20 : MUX2_X1 port map( A => Q_13_port, B => data(13), S => enable, Z => n78
                           );
   U21 : MUX2_X1 port map( A => Q_12_port, B => data(12), S => enable, Z => n77
                           );
   U22 : MUX2_X1 port map( A => Q_11_port, B => data(11), S => enable, Z => n76
                           );
   U23 : MUX2_X1 port map( A => Q_10_port, B => data(10), S => enable, Z => n75
                           );
   U24 : MUX2_X1 port map( A => Q_9_port, B => data(9), S => enable, Z => n74);
   U25 : MUX2_X1 port map( A => Q_8_port, B => data(8), S => enable, Z => n73);
   U26 : MUX2_X1 port map( A => Q_7_port, B => data(7), S => enable, Z => n72);
   U27 : MUX2_X1 port map( A => Q_6_port, B => data(6), S => enable, Z => n71);
   U28 : MUX2_X1 port map( A => Q_5_port, B => data(5), S => enable, Z => n70);
   U29 : MUX2_X1 port map( A => Q_4_port, B => data(4), S => enable, Z => n69);
   U30 : MUX2_X1 port map( A => Q_3_port, B => data(3), S => enable, Z => n68);
   U31 : MUX2_X1 port map( A => Q_2_port, B => data(2), S => enable, Z => n67);
   U32 : MUX2_X1 port map( A => Q_1_port, B => data(1), S => enable, Z => n66);
   U33 : MUX2_X1 port map( A => Q_0_port, B => data(0), S => enable, Z => n65);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity SIG_EXT_BITS32 is

   port( EXT_UNSIGNED, EXT_FOR_J : in std_logic;  S_IN : in std_logic_vector 
         (31 downto 0);  S_OUT : out std_logic_vector (31 downto 0));

end SIG_EXT_BITS32;

architecture SYN_BEHAVIOR of SIG_EXT_BITS32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal S_OUT_26_port, S_OUT_25_port, S_OUT_24_port, S_OUT_23_port, 
      S_OUT_22_port, S_OUT_21_port, S_OUT_20_port, S_OUT_19_port, S_OUT_18_port
      , S_OUT_17_port, S_OUT_16_port, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, 
      n11, n12, n13, n14 : std_logic;

begin
   S_OUT <= ( S_OUT_26_port, S_OUT_26_port, S_OUT_26_port, S_OUT_26_port, 
      S_OUT_26_port, S_OUT_26_port, S_OUT_25_port, S_OUT_24_port, S_OUT_23_port
      , S_OUT_22_port, S_OUT_21_port, S_OUT_20_port, S_OUT_19_port, 
      S_OUT_18_port, S_OUT_17_port, S_OUT_16_port, S_IN(15), S_IN(14), S_IN(13)
      , S_IN(12), S_IN(11), S_IN(10), S_IN(9), S_IN(8), S_IN(7), S_IN(6), 
      S_IN(5), S_IN(4), S_IN(3), S_IN(2), S_IN(1), S_IN(0) );
   
   U2 : NAND2_X1 port map( A1 => n1, A2 => n2, ZN => S_OUT_26_port);
   U3 : NAND3_X1 port map( A1 => EXT_FOR_J, A2 => n3, A3 => S_IN(25), ZN => n2)
                           ;
   U4 : OAI21_X1 port map( B1 => n4, B2 => n5, A => n1, ZN => S_OUT_25_port);
   U5 : INV_X1 port map( A => S_IN(25), ZN => n5);
   U6 : NAND2_X1 port map( A1 => n1, A2 => n6, ZN => S_OUT_24_port);
   U7 : NAND2_X1 port map( A1 => S_IN(24), A2 => EXT_FOR_J, ZN => n6);
   U8 : NAND2_X1 port map( A1 => n1, A2 => n7, ZN => S_OUT_23_port);
   U9 : NAND2_X1 port map( A1 => S_IN(23), A2 => EXT_FOR_J, ZN => n7);
   U10 : NAND2_X1 port map( A1 => n1, A2 => n8, ZN => S_OUT_22_port);
   U11 : NAND2_X1 port map( A1 => S_IN(22), A2 => EXT_FOR_J, ZN => n8);
   U12 : NAND2_X1 port map( A1 => n1, A2 => n9, ZN => S_OUT_21_port);
   U13 : NAND2_X1 port map( A1 => S_IN(21), A2 => EXT_FOR_J, ZN => n9);
   U14 : NAND2_X1 port map( A1 => n1, A2 => n10, ZN => S_OUT_20_port);
   U15 : NAND2_X1 port map( A1 => S_IN(20), A2 => EXT_FOR_J, ZN => n10);
   U16 : NAND2_X1 port map( A1 => n1, A2 => n11, ZN => S_OUT_19_port);
   U17 : NAND2_X1 port map( A1 => S_IN(19), A2 => EXT_FOR_J, ZN => n11);
   U18 : NAND2_X1 port map( A1 => n1, A2 => n12, ZN => S_OUT_18_port);
   U19 : NAND2_X1 port map( A1 => S_IN(18), A2 => EXT_FOR_J, ZN => n12);
   U20 : NAND2_X1 port map( A1 => n1, A2 => n13, ZN => S_OUT_17_port);
   U21 : NAND2_X1 port map( A1 => S_IN(17), A2 => EXT_FOR_J, ZN => n13);
   U22 : NAND2_X1 port map( A1 => n1, A2 => n14, ZN => S_OUT_16_port);
   U23 : NAND2_X1 port map( A1 => S_IN(16), A2 => EXT_FOR_J, ZN => n14);
   U24 : NAND3_X1 port map( A1 => n4, A2 => n3, A3 => S_IN(15), ZN => n1);
   U25 : INV_X1 port map( A => EXT_UNSIGNED, ZN => n3);
   U26 : INV_X1 port map( A => EXT_FOR_J, ZN => n4);

end SYN_BEHAVIOR;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity register_file_NBIT32_row32 is

   port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
         ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
         std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector (31
         downto 0));

end register_file_NBIT32_row32;

architecture SYN_A of register_file_NBIT32_row32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X2
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X4
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal REGISTERS_0_31_port, REGISTERS_0_30_port, REGISTERS_0_29_port, 
      REGISTERS_0_28_port, REGISTERS_0_27_port, REGISTERS_0_26_port, 
      REGISTERS_0_25_port, REGISTERS_0_24_port, REGISTERS_0_23_port, 
      REGISTERS_0_22_port, REGISTERS_0_21_port, REGISTERS_0_20_port, 
      REGISTERS_0_19_port, REGISTERS_0_18_port, REGISTERS_0_17_port, 
      REGISTERS_0_16_port, REGISTERS_0_15_port, REGISTERS_0_14_port, 
      REGISTERS_0_13_port, REGISTERS_0_12_port, REGISTERS_0_11_port, 
      REGISTERS_0_10_port, REGISTERS_0_9_port, REGISTERS_0_8_port, 
      REGISTERS_0_7_port, REGISTERS_0_6_port, REGISTERS_0_5_port, 
      REGISTERS_0_4_port, REGISTERS_0_3_port, REGISTERS_0_2_port, 
      REGISTERS_0_1_port, REGISTERS_0_0_port, REGISTERS_1_31_port, 
      REGISTERS_1_30_port, REGISTERS_1_29_port, REGISTERS_1_28_port, 
      REGISTERS_1_27_port, REGISTERS_1_26_port, REGISTERS_1_25_port, 
      REGISTERS_1_24_port, REGISTERS_1_23_port, REGISTERS_1_22_port, 
      REGISTERS_1_21_port, REGISTERS_1_20_port, REGISTERS_1_19_port, 
      REGISTERS_1_18_port, REGISTERS_1_17_port, REGISTERS_1_16_port, 
      REGISTERS_1_15_port, REGISTERS_1_14_port, REGISTERS_1_13_port, 
      REGISTERS_1_12_port, REGISTERS_1_11_port, REGISTERS_1_10_port, 
      REGISTERS_1_9_port, REGISTERS_1_8_port, REGISTERS_1_7_port, 
      REGISTERS_1_6_port, REGISTERS_1_5_port, REGISTERS_1_4_port, 
      REGISTERS_1_3_port, REGISTERS_1_2_port, REGISTERS_1_1_port, 
      REGISTERS_1_0_port, REGISTERS_2_31_port, REGISTERS_2_30_port, 
      REGISTERS_2_29_port, REGISTERS_2_28_port, REGISTERS_2_27_port, 
      REGISTERS_2_26_port, REGISTERS_2_25_port, REGISTERS_2_24_port, 
      REGISTERS_2_23_port, REGISTERS_2_22_port, REGISTERS_2_21_port, 
      REGISTERS_2_20_port, REGISTERS_2_19_port, REGISTERS_2_18_port, 
      REGISTERS_2_17_port, REGISTERS_2_16_port, REGISTERS_2_15_port, 
      REGISTERS_2_14_port, REGISTERS_2_13_port, REGISTERS_2_12_port, 
      REGISTERS_2_11_port, REGISTERS_2_10_port, REGISTERS_2_9_port, 
      REGISTERS_2_8_port, REGISTERS_2_7_port, REGISTERS_2_6_port, 
      REGISTERS_2_5_port, REGISTERS_2_4_port, REGISTERS_2_3_port, 
      REGISTERS_2_2_port, REGISTERS_2_1_port, REGISTERS_2_0_port, 
      REGISTERS_3_31_port, REGISTERS_3_30_port, REGISTERS_3_29_port, 
      REGISTERS_3_28_port, REGISTERS_3_27_port, REGISTERS_3_26_port, 
      REGISTERS_3_25_port, REGISTERS_3_24_port, REGISTERS_3_23_port, 
      REGISTERS_3_22_port, REGISTERS_3_21_port, REGISTERS_3_20_port, 
      REGISTERS_3_19_port, REGISTERS_3_18_port, REGISTERS_3_17_port, 
      REGISTERS_3_16_port, REGISTERS_3_15_port, REGISTERS_3_14_port, 
      REGISTERS_3_13_port, REGISTERS_3_12_port, REGISTERS_3_11_port, 
      REGISTERS_3_10_port, REGISTERS_3_9_port, REGISTERS_3_8_port, 
      REGISTERS_3_7_port, REGISTERS_3_6_port, REGISTERS_3_5_port, 
      REGISTERS_3_4_port, REGISTERS_3_3_port, REGISTERS_3_2_port, 
      REGISTERS_3_1_port, REGISTERS_3_0_port, REGISTERS_4_31_port, 
      REGISTERS_4_30_port, REGISTERS_4_29_port, REGISTERS_4_28_port, 
      REGISTERS_4_27_port, REGISTERS_4_26_port, REGISTERS_4_25_port, 
      REGISTERS_4_24_port, REGISTERS_4_23_port, REGISTERS_4_22_port, 
      REGISTERS_4_21_port, REGISTERS_4_20_port, REGISTERS_4_19_port, 
      REGISTERS_4_18_port, REGISTERS_4_17_port, REGISTERS_4_16_port, 
      REGISTERS_4_15_port, REGISTERS_4_14_port, REGISTERS_4_13_port, 
      REGISTERS_4_12_port, REGISTERS_4_11_port, REGISTERS_4_10_port, 
      REGISTERS_4_9_port, REGISTERS_4_8_port, REGISTERS_4_7_port, 
      REGISTERS_4_6_port, REGISTERS_4_5_port, REGISTERS_4_4_port, 
      REGISTERS_4_3_port, REGISTERS_4_2_port, REGISTERS_4_1_port, 
      REGISTERS_4_0_port, REGISTERS_5_31_port, REGISTERS_5_30_port, 
      REGISTERS_5_29_port, REGISTERS_5_28_port, REGISTERS_5_27_port, 
      REGISTERS_5_26_port, REGISTERS_5_25_port, REGISTERS_5_24_port, 
      REGISTERS_5_23_port, REGISTERS_5_22_port, REGISTERS_5_21_port, 
      REGISTERS_5_20_port, REGISTERS_5_19_port, REGISTERS_5_18_port, 
      REGISTERS_5_17_port, REGISTERS_5_16_port, REGISTERS_5_15_port, 
      REGISTERS_5_14_port, REGISTERS_5_13_port, REGISTERS_5_12_port, 
      REGISTERS_5_11_port, REGISTERS_5_10_port, REGISTERS_5_9_port, 
      REGISTERS_5_8_port, REGISTERS_5_7_port, REGISTERS_5_6_port, 
      REGISTERS_5_5_port, REGISTERS_5_4_port, REGISTERS_5_3_port, 
      REGISTERS_5_2_port, REGISTERS_5_1_port, REGISTERS_5_0_port, 
      REGISTERS_6_31_port, REGISTERS_6_30_port, REGISTERS_6_29_port, 
      REGISTERS_6_28_port, REGISTERS_6_27_port, REGISTERS_6_26_port, 
      REGISTERS_6_25_port, REGISTERS_6_24_port, REGISTERS_6_23_port, 
      REGISTERS_6_22_port, REGISTERS_6_21_port, REGISTERS_6_20_port, 
      REGISTERS_6_19_port, REGISTERS_6_18_port, REGISTERS_6_17_port, 
      REGISTERS_6_16_port, REGISTERS_6_15_port, REGISTERS_6_14_port, 
      REGISTERS_6_13_port, REGISTERS_6_12_port, REGISTERS_6_11_port, 
      REGISTERS_6_10_port, REGISTERS_6_9_port, REGISTERS_6_8_port, 
      REGISTERS_6_7_port, REGISTERS_6_6_port, REGISTERS_6_5_port, 
      REGISTERS_6_4_port, REGISTERS_6_3_port, REGISTERS_6_2_port, 
      REGISTERS_6_1_port, REGISTERS_6_0_port, REGISTERS_7_31_port, 
      REGISTERS_7_30_port, REGISTERS_7_29_port, REGISTERS_7_28_port, 
      REGISTERS_7_27_port, REGISTERS_7_26_port, REGISTERS_7_25_port, 
      REGISTERS_7_24_port, REGISTERS_7_23_port, REGISTERS_7_22_port, 
      REGISTERS_7_21_port, REGISTERS_7_20_port, REGISTERS_7_19_port, 
      REGISTERS_7_18_port, REGISTERS_7_17_port, REGISTERS_7_16_port, 
      REGISTERS_7_15_port, REGISTERS_7_14_port, REGISTERS_7_13_port, 
      REGISTERS_7_12_port, REGISTERS_7_11_port, REGISTERS_7_10_port, 
      REGISTERS_7_9_port, REGISTERS_7_8_port, REGISTERS_7_7_port, 
      REGISTERS_7_6_port, REGISTERS_7_5_port, REGISTERS_7_4_port, 
      REGISTERS_7_3_port, REGISTERS_7_2_port, REGISTERS_7_1_port, 
      REGISTERS_7_0_port, REGISTERS_8_31_port, REGISTERS_8_30_port, 
      REGISTERS_8_29_port, REGISTERS_8_28_port, REGISTERS_8_27_port, 
      REGISTERS_8_26_port, REGISTERS_8_25_port, REGISTERS_8_24_port, 
      REGISTERS_8_23_port, REGISTERS_8_22_port, REGISTERS_8_21_port, 
      REGISTERS_8_20_port, REGISTERS_8_19_port, REGISTERS_8_18_port, 
      REGISTERS_8_17_port, REGISTERS_8_16_port, REGISTERS_8_15_port, 
      REGISTERS_8_14_port, REGISTERS_8_13_port, REGISTERS_8_12_port, 
      REGISTERS_8_11_port, REGISTERS_8_10_port, REGISTERS_8_9_port, 
      REGISTERS_8_8_port, REGISTERS_8_7_port, REGISTERS_8_6_port, 
      REGISTERS_8_5_port, REGISTERS_8_4_port, REGISTERS_8_3_port, 
      REGISTERS_8_2_port, REGISTERS_8_1_port, REGISTERS_8_0_port, 
      REGISTERS_9_31_port, REGISTERS_9_30_port, REGISTERS_9_29_port, 
      REGISTERS_9_28_port, REGISTERS_9_27_port, REGISTERS_9_26_port, 
      REGISTERS_9_25_port, REGISTERS_9_24_port, REGISTERS_9_23_port, 
      REGISTERS_9_22_port, REGISTERS_9_21_port, REGISTERS_9_20_port, 
      REGISTERS_9_19_port, REGISTERS_9_18_port, REGISTERS_9_17_port, 
      REGISTERS_9_16_port, REGISTERS_9_15_port, REGISTERS_9_14_port, 
      REGISTERS_9_13_port, REGISTERS_9_12_port, REGISTERS_9_11_port, 
      REGISTERS_9_10_port, REGISTERS_9_9_port, REGISTERS_9_8_port, 
      REGISTERS_9_7_port, REGISTERS_9_6_port, REGISTERS_9_5_port, 
      REGISTERS_9_4_port, REGISTERS_9_3_port, REGISTERS_9_2_port, 
      REGISTERS_9_1_port, REGISTERS_9_0_port, REGISTERS_10_31_port, 
      REGISTERS_10_30_port, REGISTERS_10_29_port, REGISTERS_10_28_port, 
      REGISTERS_10_27_port, REGISTERS_10_26_port, REGISTERS_10_25_port, 
      REGISTERS_10_24_port, REGISTERS_10_23_port, REGISTERS_10_22_port, 
      REGISTERS_10_21_port, REGISTERS_10_20_port, REGISTERS_10_19_port, 
      REGISTERS_10_18_port, REGISTERS_10_17_port, REGISTERS_10_16_port, 
      REGISTERS_10_15_port, REGISTERS_10_14_port, REGISTERS_10_13_port, 
      REGISTERS_10_12_port, REGISTERS_10_11_port, REGISTERS_10_10_port, 
      REGISTERS_10_9_port, REGISTERS_10_8_port, REGISTERS_10_7_port, 
      REGISTERS_10_6_port, REGISTERS_10_5_port, REGISTERS_10_4_port, 
      REGISTERS_10_3_port, REGISTERS_10_2_port, REGISTERS_10_1_port, 
      REGISTERS_10_0_port, REGISTERS_11_31_port, REGISTERS_11_30_port, 
      REGISTERS_11_29_port, REGISTERS_11_28_port, REGISTERS_11_27_port, 
      REGISTERS_11_26_port, REGISTERS_11_25_port, REGISTERS_11_24_port, 
      REGISTERS_11_23_port, REGISTERS_11_22_port, REGISTERS_11_21_port, 
      REGISTERS_11_20_port, REGISTERS_11_19_port, REGISTERS_11_18_port, 
      REGISTERS_11_17_port, REGISTERS_11_16_port, REGISTERS_11_15_port, 
      REGISTERS_11_14_port, REGISTERS_11_13_port, REGISTERS_11_12_port, 
      REGISTERS_11_11_port, REGISTERS_11_10_port, REGISTERS_11_9_port, 
      REGISTERS_11_8_port, REGISTERS_11_7_port, REGISTERS_11_6_port, 
      REGISTERS_11_5_port, REGISTERS_11_4_port, REGISTERS_11_3_port, 
      REGISTERS_11_2_port, REGISTERS_11_1_port, REGISTERS_11_0_port, 
      REGISTERS_12_31_port, REGISTERS_12_30_port, REGISTERS_12_29_port, 
      REGISTERS_12_28_port, REGISTERS_12_27_port, REGISTERS_12_26_port, 
      REGISTERS_12_25_port, REGISTERS_12_24_port, REGISTERS_12_23_port, 
      REGISTERS_12_22_port, REGISTERS_12_21_port, REGISTERS_12_20_port, 
      REGISTERS_12_19_port, REGISTERS_12_18_port, REGISTERS_12_17_port, 
      REGISTERS_12_16_port, REGISTERS_12_15_port, REGISTERS_12_14_port, 
      REGISTERS_12_13_port, REGISTERS_12_12_port, REGISTERS_12_11_port, 
      REGISTERS_12_10_port, REGISTERS_12_9_port, REGISTERS_12_8_port, 
      REGISTERS_12_7_port, REGISTERS_12_6_port, REGISTERS_12_5_port, 
      REGISTERS_12_4_port, REGISTERS_12_3_port, REGISTERS_12_2_port, 
      REGISTERS_12_1_port, REGISTERS_12_0_port, REGISTERS_13_31_port, 
      REGISTERS_13_30_port, REGISTERS_13_29_port, REGISTERS_13_28_port, 
      REGISTERS_13_27_port, REGISTERS_13_26_port, REGISTERS_13_25_port, 
      REGISTERS_13_24_port, REGISTERS_13_23_port, REGISTERS_13_22_port, 
      REGISTERS_13_21_port, REGISTERS_13_20_port, REGISTERS_13_19_port, 
      REGISTERS_13_18_port, REGISTERS_13_17_port, REGISTERS_13_16_port, 
      REGISTERS_13_15_port, REGISTERS_13_14_port, REGISTERS_13_13_port, 
      REGISTERS_13_12_port, REGISTERS_13_11_port, REGISTERS_13_10_port, 
      REGISTERS_13_9_port, REGISTERS_13_8_port, REGISTERS_13_7_port, 
      REGISTERS_13_6_port, REGISTERS_13_5_port, REGISTERS_13_4_port, 
      REGISTERS_13_3_port, REGISTERS_13_2_port, REGISTERS_13_1_port, 
      REGISTERS_13_0_port, REGISTERS_14_31_port, REGISTERS_14_30_port, 
      REGISTERS_14_29_port, REGISTERS_14_28_port, REGISTERS_14_27_port, 
      REGISTERS_14_26_port, REGISTERS_14_25_port, REGISTERS_14_24_port, 
      REGISTERS_14_23_port, REGISTERS_14_22_port, REGISTERS_14_21_port, 
      REGISTERS_14_20_port, REGISTERS_14_19_port, REGISTERS_14_18_port, 
      REGISTERS_14_17_port, REGISTERS_14_16_port, REGISTERS_14_15_port, 
      REGISTERS_14_14_port, REGISTERS_14_13_port, REGISTERS_14_12_port, 
      REGISTERS_14_11_port, REGISTERS_14_10_port, REGISTERS_14_9_port, 
      REGISTERS_14_8_port, REGISTERS_14_7_port, REGISTERS_14_6_port, 
      REGISTERS_14_5_port, REGISTERS_14_4_port, REGISTERS_14_3_port, 
      REGISTERS_14_2_port, REGISTERS_14_1_port, REGISTERS_14_0_port, 
      REGISTERS_15_31_port, REGISTERS_15_30_port, REGISTERS_15_29_port, 
      REGISTERS_15_28_port, REGISTERS_15_27_port, REGISTERS_15_26_port, 
      REGISTERS_15_25_port, REGISTERS_15_24_port, REGISTERS_15_23_port, 
      REGISTERS_15_22_port, REGISTERS_15_21_port, REGISTERS_15_20_port, 
      REGISTERS_15_19_port, REGISTERS_15_18_port, REGISTERS_15_17_port, 
      REGISTERS_15_16_port, REGISTERS_15_15_port, REGISTERS_15_14_port, 
      REGISTERS_15_13_port, REGISTERS_15_12_port, REGISTERS_15_11_port, 
      REGISTERS_15_10_port, REGISTERS_15_9_port, REGISTERS_15_8_port, 
      REGISTERS_15_7_port, REGISTERS_15_6_port, REGISTERS_15_5_port, 
      REGISTERS_15_4_port, REGISTERS_15_3_port, REGISTERS_15_2_port, 
      REGISTERS_15_1_port, REGISTERS_15_0_port, REGISTERS_16_31_port, 
      REGISTERS_16_30_port, REGISTERS_16_29_port, REGISTERS_16_28_port, 
      REGISTERS_16_27_port, REGISTERS_16_26_port, REGISTERS_16_25_port, 
      REGISTERS_16_24_port, REGISTERS_16_23_port, REGISTERS_16_22_port, 
      REGISTERS_16_21_port, REGISTERS_16_20_port, REGISTERS_16_19_port, 
      REGISTERS_16_18_port, REGISTERS_16_17_port, REGISTERS_16_16_port, 
      REGISTERS_16_15_port, REGISTERS_16_14_port, REGISTERS_16_13_port, 
      REGISTERS_16_12_port, REGISTERS_16_11_port, REGISTERS_16_10_port, 
      REGISTERS_16_9_port, REGISTERS_16_8_port, REGISTERS_16_7_port, 
      REGISTERS_16_6_port, REGISTERS_16_5_port, REGISTERS_16_4_port, 
      REGISTERS_16_3_port, REGISTERS_16_2_port, REGISTERS_16_1_port, 
      REGISTERS_16_0_port, REGISTERS_17_31_port, REGISTERS_17_30_port, 
      REGISTERS_17_29_port, REGISTERS_17_28_port, REGISTERS_17_27_port, 
      REGISTERS_17_26_port, REGISTERS_17_25_port, REGISTERS_17_24_port, 
      REGISTERS_17_23_port, REGISTERS_17_22_port, REGISTERS_17_21_port, 
      REGISTERS_17_20_port, REGISTERS_17_19_port, REGISTERS_17_18_port, 
      REGISTERS_17_17_port, REGISTERS_17_16_port, REGISTERS_17_15_port, 
      REGISTERS_17_14_port, REGISTERS_17_13_port, REGISTERS_17_12_port, 
      REGISTERS_17_11_port, REGISTERS_17_10_port, REGISTERS_17_9_port, 
      REGISTERS_17_8_port, REGISTERS_17_7_port, REGISTERS_17_6_port, 
      REGISTERS_17_5_port, REGISTERS_17_4_port, REGISTERS_17_3_port, 
      REGISTERS_17_2_port, REGISTERS_17_1_port, REGISTERS_17_0_port, 
      REGISTERS_18_31_port, REGISTERS_18_30_port, REGISTERS_18_29_port, 
      REGISTERS_18_28_port, REGISTERS_18_27_port, REGISTERS_18_26_port, 
      REGISTERS_18_25_port, REGISTERS_18_24_port, REGISTERS_18_23_port, 
      REGISTERS_18_22_port, REGISTERS_18_21_port, REGISTERS_18_20_port, 
      REGISTERS_18_19_port, REGISTERS_18_18_port, REGISTERS_18_17_port, 
      REGISTERS_18_16_port, REGISTERS_18_15_port, REGISTERS_18_14_port, 
      REGISTERS_18_13_port, REGISTERS_18_12_port, REGISTERS_18_11_port, 
      REGISTERS_18_10_port, REGISTERS_18_9_port, REGISTERS_18_8_port, 
      REGISTERS_18_7_port, REGISTERS_18_6_port, REGISTERS_18_5_port, 
      REGISTERS_18_4_port, REGISTERS_18_3_port, REGISTERS_18_2_port, 
      REGISTERS_18_1_port, REGISTERS_18_0_port, REGISTERS_19_31_port, 
      REGISTERS_19_30_port, REGISTERS_19_29_port, REGISTERS_19_28_port, 
      REGISTERS_19_27_port, REGISTERS_19_26_port, REGISTERS_19_25_port, 
      REGISTERS_19_24_port, REGISTERS_19_23_port, REGISTERS_19_22_port, 
      REGISTERS_19_21_port, REGISTERS_19_20_port, REGISTERS_19_19_port, 
      REGISTERS_19_18_port, REGISTERS_19_17_port, REGISTERS_19_16_port, 
      REGISTERS_19_15_port, REGISTERS_19_14_port, REGISTERS_19_13_port, 
      REGISTERS_19_12_port, REGISTERS_19_11_port, REGISTERS_19_10_port, 
      REGISTERS_19_9_port, REGISTERS_19_8_port, REGISTERS_19_7_port, 
      REGISTERS_19_6_port, REGISTERS_19_5_port, REGISTERS_19_4_port, 
      REGISTERS_19_3_port, REGISTERS_19_2_port, REGISTERS_19_1_port, 
      REGISTERS_19_0_port, REGISTERS_20_31_port, REGISTERS_20_30_port, 
      REGISTERS_20_29_port, REGISTERS_20_28_port, REGISTERS_20_27_port, 
      REGISTERS_20_26_port, REGISTERS_20_25_port, REGISTERS_20_24_port, 
      REGISTERS_20_23_port, REGISTERS_20_22_port, REGISTERS_20_21_port, 
      REGISTERS_20_20_port, REGISTERS_20_19_port, REGISTERS_20_18_port, 
      REGISTERS_20_17_port, REGISTERS_20_16_port, REGISTERS_20_15_port, 
      REGISTERS_20_14_port, REGISTERS_20_13_port, REGISTERS_20_12_port, 
      REGISTERS_20_11_port, REGISTERS_20_10_port, REGISTERS_20_9_port, 
      REGISTERS_20_8_port, REGISTERS_20_7_port, REGISTERS_20_6_port, 
      REGISTERS_20_5_port, REGISTERS_20_4_port, REGISTERS_20_3_port, 
      REGISTERS_20_2_port, REGISTERS_20_1_port, REGISTERS_20_0_port, 
      REGISTERS_21_31_port, REGISTERS_21_30_port, REGISTERS_21_29_port, 
      REGISTERS_21_28_port, REGISTERS_21_27_port, REGISTERS_21_26_port, 
      REGISTERS_21_25_port, REGISTERS_21_24_port, REGISTERS_21_23_port, 
      REGISTERS_21_22_port, REGISTERS_21_21_port, REGISTERS_21_20_port, 
      REGISTERS_21_19_port, REGISTERS_21_18_port, REGISTERS_21_17_port, 
      REGISTERS_21_16_port, REGISTERS_21_15_port, REGISTERS_21_14_port, 
      REGISTERS_21_13_port, REGISTERS_21_12_port, REGISTERS_21_11_port, 
      REGISTERS_21_10_port, REGISTERS_21_9_port, REGISTERS_21_8_port, 
      REGISTERS_21_7_port, REGISTERS_21_6_port, REGISTERS_21_5_port, 
      REGISTERS_21_4_port, REGISTERS_21_3_port, REGISTERS_21_2_port, 
      REGISTERS_21_1_port, REGISTERS_21_0_port, REGISTERS_22_31_port, 
      REGISTERS_22_30_port, REGISTERS_22_29_port, REGISTERS_22_28_port, 
      REGISTERS_22_27_port, REGISTERS_22_26_port, REGISTERS_22_25_port, 
      REGISTERS_22_24_port, REGISTERS_22_23_port, REGISTERS_22_22_port, 
      REGISTERS_22_21_port, REGISTERS_22_20_port, REGISTERS_22_19_port, 
      REGISTERS_22_18_port, REGISTERS_22_17_port, REGISTERS_22_16_port, 
      REGISTERS_22_15_port, REGISTERS_22_14_port, REGISTERS_22_13_port, 
      REGISTERS_22_12_port, REGISTERS_22_11_port, REGISTERS_22_10_port, 
      REGISTERS_22_9_port, REGISTERS_22_8_port, REGISTERS_22_7_port, 
      REGISTERS_22_6_port, REGISTERS_22_5_port, REGISTERS_22_4_port, 
      REGISTERS_22_3_port, REGISTERS_22_2_port, REGISTERS_22_1_port, 
      REGISTERS_22_0_port, REGISTERS_23_31_port, REGISTERS_23_30_port, 
      REGISTERS_23_29_port, REGISTERS_23_28_port, REGISTERS_23_27_port, 
      REGISTERS_23_26_port, REGISTERS_23_25_port, REGISTERS_23_24_port, 
      REGISTERS_23_23_port, REGISTERS_23_22_port, REGISTERS_23_21_port, 
      REGISTERS_23_20_port, REGISTERS_23_19_port, REGISTERS_23_18_port, 
      REGISTERS_23_17_port, REGISTERS_23_16_port, REGISTERS_23_15_port, 
      REGISTERS_23_14_port, REGISTERS_23_13_port, REGISTERS_23_12_port, 
      REGISTERS_23_11_port, REGISTERS_23_10_port, REGISTERS_23_9_port, 
      REGISTERS_23_8_port, REGISTERS_23_7_port, REGISTERS_23_6_port, 
      REGISTERS_23_5_port, REGISTERS_23_4_port, REGISTERS_23_3_port, 
      REGISTERS_23_2_port, REGISTERS_23_1_port, REGISTERS_23_0_port, 
      REGISTERS_24_31_port, REGISTERS_24_30_port, REGISTERS_24_29_port, 
      REGISTERS_24_28_port, REGISTERS_24_27_port, REGISTERS_24_26_port, 
      REGISTERS_24_25_port, REGISTERS_24_24_port, REGISTERS_24_23_port, 
      REGISTERS_24_22_port, REGISTERS_24_21_port, REGISTERS_24_20_port, 
      REGISTERS_24_19_port, REGISTERS_24_18_port, REGISTERS_24_17_port, 
      REGISTERS_24_16_port, REGISTERS_24_15_port, REGISTERS_24_14_port, 
      REGISTERS_24_13_port, REGISTERS_24_12_port, REGISTERS_24_11_port, 
      REGISTERS_24_10_port, REGISTERS_24_9_port, REGISTERS_24_8_port, 
      REGISTERS_24_7_port, REGISTERS_24_6_port, REGISTERS_24_5_port, 
      REGISTERS_24_4_port, REGISTERS_24_3_port, REGISTERS_24_2_port, 
      REGISTERS_24_1_port, REGISTERS_24_0_port, REGISTERS_25_31_port, 
      REGISTERS_25_30_port, REGISTERS_25_29_port, REGISTERS_25_28_port, 
      REGISTERS_25_27_port, REGISTERS_25_26_port, REGISTERS_25_25_port, 
      REGISTERS_25_24_port, REGISTERS_25_23_port, REGISTERS_25_22_port, 
      REGISTERS_25_21_port, REGISTERS_25_20_port, REGISTERS_25_19_port, 
      REGISTERS_25_18_port, REGISTERS_25_17_port, REGISTERS_25_16_port, 
      REGISTERS_25_15_port, REGISTERS_25_14_port, REGISTERS_25_13_port, 
      REGISTERS_25_12_port, REGISTERS_25_11_port, REGISTERS_25_10_port, 
      REGISTERS_25_9_port, REGISTERS_25_8_port, REGISTERS_25_7_port, 
      REGISTERS_25_6_port, REGISTERS_25_5_port, REGISTERS_25_4_port, 
      REGISTERS_25_3_port, REGISTERS_25_2_port, REGISTERS_25_1_port, 
      REGISTERS_25_0_port, REGISTERS_26_31_port, REGISTERS_26_30_port, 
      REGISTERS_26_29_port, REGISTERS_26_28_port, REGISTERS_26_27_port, 
      REGISTERS_26_26_port, REGISTERS_26_25_port, REGISTERS_26_24_port, 
      REGISTERS_26_23_port, REGISTERS_26_22_port, REGISTERS_26_21_port, 
      REGISTERS_26_20_port, REGISTERS_26_19_port, REGISTERS_26_18_port, 
      REGISTERS_26_17_port, REGISTERS_26_16_port, REGISTERS_26_15_port, 
      REGISTERS_26_14_port, REGISTERS_26_13_port, REGISTERS_26_12_port, 
      REGISTERS_26_11_port, REGISTERS_26_10_port, REGISTERS_26_9_port, 
      REGISTERS_26_8_port, REGISTERS_26_7_port, REGISTERS_26_6_port, 
      REGISTERS_26_5_port, REGISTERS_26_4_port, REGISTERS_26_3_port, 
      REGISTERS_26_2_port, REGISTERS_26_1_port, REGISTERS_26_0_port, 
      REGISTERS_27_31_port, REGISTERS_27_30_port, REGISTERS_27_29_port, 
      REGISTERS_27_28_port, REGISTERS_27_27_port, REGISTERS_27_26_port, 
      REGISTERS_27_25_port, REGISTERS_27_24_port, REGISTERS_27_23_port, 
      REGISTERS_27_22_port, REGISTERS_27_21_port, REGISTERS_27_20_port, 
      REGISTERS_27_19_port, REGISTERS_27_18_port, REGISTERS_27_17_port, 
      REGISTERS_27_16_port, REGISTERS_27_15_port, REGISTERS_27_14_port, 
      REGISTERS_27_13_port, REGISTERS_27_12_port, REGISTERS_27_11_port, 
      REGISTERS_27_10_port, REGISTERS_27_9_port, REGISTERS_27_8_port, 
      REGISTERS_27_7_port, REGISTERS_27_6_port, REGISTERS_27_5_port, 
      REGISTERS_27_4_port, REGISTERS_27_3_port, REGISTERS_27_2_port, 
      REGISTERS_27_1_port, REGISTERS_27_0_port, REGISTERS_28_31_port, 
      REGISTERS_28_30_port, REGISTERS_28_29_port, REGISTERS_28_28_port, 
      REGISTERS_28_27_port, REGISTERS_28_26_port, REGISTERS_28_25_port, 
      REGISTERS_28_24_port, REGISTERS_28_23_port, REGISTERS_28_22_port, 
      REGISTERS_28_21_port, REGISTERS_28_20_port, REGISTERS_28_19_port, 
      REGISTERS_28_18_port, REGISTERS_28_17_port, REGISTERS_28_16_port, 
      REGISTERS_28_15_port, REGISTERS_28_14_port, REGISTERS_28_13_port, 
      REGISTERS_28_12_port, REGISTERS_28_11_port, REGISTERS_28_10_port, 
      REGISTERS_28_9_port, REGISTERS_28_8_port, REGISTERS_28_7_port, 
      REGISTERS_28_6_port, REGISTERS_28_5_port, REGISTERS_28_4_port, 
      REGISTERS_28_3_port, REGISTERS_28_2_port, REGISTERS_28_1_port, 
      REGISTERS_28_0_port, REGISTERS_29_31_port, REGISTERS_29_30_port, 
      REGISTERS_29_29_port, REGISTERS_29_28_port, REGISTERS_29_27_port, 
      REGISTERS_29_26_port, REGISTERS_29_25_port, REGISTERS_29_24_port, 
      REGISTERS_29_23_port, REGISTERS_29_22_port, REGISTERS_29_21_port, 
      REGISTERS_29_20_port, REGISTERS_29_19_port, REGISTERS_29_18_port, 
      REGISTERS_29_17_port, REGISTERS_29_16_port, REGISTERS_29_15_port, 
      REGISTERS_29_14_port, REGISTERS_29_13_port, REGISTERS_29_12_port, 
      REGISTERS_29_11_port, REGISTERS_29_10_port, REGISTERS_29_9_port, 
      REGISTERS_29_8_port, REGISTERS_29_7_port, REGISTERS_29_6_port, 
      REGISTERS_29_5_port, REGISTERS_29_4_port, REGISTERS_29_3_port, 
      REGISTERS_29_2_port, REGISTERS_29_1_port, REGISTERS_29_0_port, 
      REGISTERS_30_31_port, REGISTERS_30_30_port, REGISTERS_30_29_port, 
      REGISTERS_30_28_port, REGISTERS_30_27_port, REGISTERS_30_26_port, 
      REGISTERS_30_25_port, REGISTERS_30_24_port, REGISTERS_30_23_port, 
      REGISTERS_30_22_port, REGISTERS_30_21_port, REGISTERS_30_20_port, 
      REGISTERS_30_19_port, REGISTERS_30_18_port, REGISTERS_30_17_port, 
      REGISTERS_30_16_port, REGISTERS_30_15_port, REGISTERS_30_14_port, 
      REGISTERS_30_13_port, REGISTERS_30_12_port, REGISTERS_30_11_port, 
      REGISTERS_30_10_port, REGISTERS_30_9_port, REGISTERS_30_8_port, 
      REGISTERS_30_7_port, REGISTERS_30_6_port, REGISTERS_30_5_port, 
      REGISTERS_30_4_port, REGISTERS_30_3_port, REGISTERS_30_2_port, 
      REGISTERS_30_1_port, REGISTERS_30_0_port, REGISTERS_31_31_port, 
      REGISTERS_31_30_port, REGISTERS_31_29_port, REGISTERS_31_28_port, 
      REGISTERS_31_27_port, REGISTERS_31_26_port, REGISTERS_31_25_port, 
      REGISTERS_31_24_port, REGISTERS_31_23_port, REGISTERS_31_22_port, 
      REGISTERS_31_21_port, REGISTERS_31_20_port, REGISTERS_31_19_port, 
      REGISTERS_31_18_port, REGISTERS_31_17_port, REGISTERS_31_16_port, 
      REGISTERS_31_15_port, REGISTERS_31_14_port, REGISTERS_31_13_port, 
      REGISTERS_31_12_port, REGISTERS_31_11_port, REGISTERS_31_10_port, 
      REGISTERS_31_9_port, REGISTERS_31_8_port, REGISTERS_31_7_port, 
      REGISTERS_31_6_port, REGISTERS_31_5_port, REGISTERS_31_4_port, 
      REGISTERS_31_3_port, REGISTERS_31_2_port, REGISTERS_31_1_port, 
      REGISTERS_31_0_port, N2419, N2421, N2423, N2425, N2427, N2429, N2431, 
      N2433, N2435, N2437, N2439, N2441, N2443, N2445, N2447, N2449, N2451, 
      N2453, N2455, N2457, N2459, N2461, N2463, N2465, N2467, N2469, N2471, 
      N2473, N2475, N2477, N2479, N2480, N2481, N2483, N2485, N2487, N2489, 
      N2491, N2493, N2495, N2497, N2499, N2501, N2503, N2505, N2507, N2509, 
      N2511, N2513, N2515, N2517, N2519, N2521, N2523, N2525, N2527, N2529, 
      N2531, N2533, N2535, N2537, N2539, N2541, N2543, N2544, N2545, N2608, 
      N2672, N2736, N2800, N2864, N2928, N2992, N3056, N3120, N3184, N3248, 
      N3312, N3376, N3440, N3504, N3568, N3632, N3696, N3760, N3824, N3888, 
      N3952, N4016, N4080, N4144, N4208, N4272, N4336, N4400, N4464, N4528, 
      N4531, N4533, N4535, N4537, N4539, N4541, N4543, N4545, N4547, N4549, 
      N4551, N4553, N4555, N4557, N4559, N4561, N4563, N4565, N4567, N4569, 
      N4571, N4573, N4575, N4577, N4579, N4581, N4583, N4585, N4587, N4589, 
      N4591, N4592, N4593, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, 
      n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27
      , n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, 
      n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56
      , n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, 
      n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85
      , n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, 
      n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, 
      n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, 
      n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, 
      n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, 
      n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, 
      n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, 
      n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, 
      n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, 
      n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, 
      n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, 
      n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, 
      n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, 
      n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, 
      n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, 
      n268, n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, 
      n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, 
      n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, 
      n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, 
      n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327, 
      n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, 
      n340, n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, 
      n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, 
      n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, 
      n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, 
      n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, 
      n400, n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, 
      n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, 
      n424, n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, 
      n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, 
      n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, 
      n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, 
      n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, 
      n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, 
      n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, 
      n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519, 
      n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, 
      n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543, 
      n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, 
      n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, 
      n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, 
      n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591, 
      n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, 
      n604, n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, 
      n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, 
      n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, 
      n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, 
      n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, 
      n664, n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, 
      n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, 
      n688, n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, 
      n700, n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, 
      n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, 
      n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, 
      n736, n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, 
      n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, 
      n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, 
      n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, 
      n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, 
      n796, n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, 
      n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, 
      n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, 
      n832, n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, 
      n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, 
      n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, 
      n868, n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, 
      n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, 
      n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, 
      n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, 
      n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, 
      n928, n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, 
      n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, 
      n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, 
      n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, 
      n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, 
      n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, 
      n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, 
      n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, 
      n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, 
      n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, 
      n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, 
      n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, 
      n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, 
      n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, 
      n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, 
      n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, 
      n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, 
      n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, 
      n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, 
      n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, 
      n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, 
      n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, 
      n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, 
      n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, 
      n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, 
      n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, 
      n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, 
      n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, 
      n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, 
      n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, 
      n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, 
      n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, 
      n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, 
      n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, 
      n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, 
      n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, 
      n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, 
      n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, 
      n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, 
      n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, 
      n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, 
      n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, 
      n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, 
      n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, 
      n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, 
      n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, 
      n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, 
      n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, 
      n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, 
      n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, 
      n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, 
      n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, 
      n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, 
      n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, 
      n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, 
      n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, 
      n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, 
      n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, 
      n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, 
      n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, 
      n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, 
      n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, 
      n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, 
      n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, 
      n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, 
      n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, 
      n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, 
      n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, 
      n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, 
      n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, 
      n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, 
      n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, 
      n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, 
      n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, 
      n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, 
      n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, 
      n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, 
      n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, 
      n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, 
      n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, 
      n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, 
      n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, 
      n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, 
      n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778 : std_logic
      ;

begin
   
   REGISTERS_reg_0_31_inst : DLH_X1 port map( G => N4592, D => N4593, Q => 
                           REGISTERS_0_31_port);
   REGISTERS_reg_0_30_inst : DLH_X1 port map( G => N4592, D => N4591, Q => 
                           REGISTERS_0_30_port);
   REGISTERS_reg_0_29_inst : DLH_X1 port map( G => N4592, D => N4589, Q => 
                           REGISTERS_0_29_port);
   REGISTERS_reg_0_28_inst : DLH_X1 port map( G => N4592, D => N4587, Q => 
                           REGISTERS_0_28_port);
   REGISTERS_reg_0_27_inst : DLH_X1 port map( G => N4592, D => N4585, Q => 
                           REGISTERS_0_27_port);
   REGISTERS_reg_0_26_inst : DLH_X1 port map( G => N4592, D => N4583, Q => 
                           REGISTERS_0_26_port);
   REGISTERS_reg_0_25_inst : DLH_X1 port map( G => N4592, D => N4581, Q => 
                           REGISTERS_0_25_port);
   REGISTERS_reg_0_24_inst : DLH_X1 port map( G => N4592, D => N4579, Q => 
                           REGISTERS_0_24_port);
   REGISTERS_reg_0_23_inst : DLH_X1 port map( G => N4592, D => N4577, Q => 
                           REGISTERS_0_23_port);
   REGISTERS_reg_0_22_inst : DLH_X1 port map( G => N4592, D => N4575, Q => 
                           REGISTERS_0_22_port);
   REGISTERS_reg_0_21_inst : DLH_X1 port map( G => N4592, D => N4573, Q => 
                           REGISTERS_0_21_port);
   REGISTERS_reg_0_20_inst : DLH_X1 port map( G => N4592, D => N4571, Q => 
                           REGISTERS_0_20_port);
   REGISTERS_reg_0_19_inst : DLH_X1 port map( G => N4592, D => N4569, Q => 
                           REGISTERS_0_19_port);
   REGISTERS_reg_0_18_inst : DLH_X1 port map( G => N4592, D => N4567, Q => 
                           REGISTERS_0_18_port);
   REGISTERS_reg_0_17_inst : DLH_X1 port map( G => N4592, D => N4565, Q => 
                           REGISTERS_0_17_port);
   REGISTERS_reg_0_16_inst : DLH_X1 port map( G => N4592, D => N4563, Q => 
                           REGISTERS_0_16_port);
   REGISTERS_reg_0_15_inst : DLH_X1 port map( G => N4592, D => N4561, Q => 
                           REGISTERS_0_15_port);
   REGISTERS_reg_0_14_inst : DLH_X1 port map( G => N4592, D => N4559, Q => 
                           REGISTERS_0_14_port);
   REGISTERS_reg_0_13_inst : DLH_X1 port map( G => N4592, D => N4557, Q => 
                           REGISTERS_0_13_port);
   REGISTERS_reg_0_12_inst : DLH_X1 port map( G => N4592, D => N4555, Q => 
                           REGISTERS_0_12_port);
   REGISTERS_reg_0_11_inst : DLH_X1 port map( G => N4592, D => N4553, Q => 
                           REGISTERS_0_11_port);
   REGISTERS_reg_0_10_inst : DLH_X1 port map( G => N4592, D => N4551, Q => 
                           REGISTERS_0_10_port);
   REGISTERS_reg_0_9_inst : DLH_X1 port map( G => N4592, D => N4549, Q => 
                           REGISTERS_0_9_port);
   REGISTERS_reg_0_8_inst : DLH_X1 port map( G => N4592, D => N4547, Q => 
                           REGISTERS_0_8_port);
   REGISTERS_reg_0_7_inst : DLH_X1 port map( G => N4592, D => N4545, Q => 
                           REGISTERS_0_7_port);
   REGISTERS_reg_0_6_inst : DLH_X1 port map( G => N4592, D => N4543, Q => 
                           REGISTERS_0_6_port);
   REGISTERS_reg_0_5_inst : DLH_X1 port map( G => N4592, D => N4541, Q => 
                           REGISTERS_0_5_port);
   REGISTERS_reg_0_4_inst : DLH_X1 port map( G => N4592, D => N4539, Q => 
                           REGISTERS_0_4_port);
   REGISTERS_reg_0_3_inst : DLH_X1 port map( G => N4592, D => N4537, Q => 
                           REGISTERS_0_3_port);
   REGISTERS_reg_0_2_inst : DLH_X1 port map( G => N4592, D => N4535, Q => 
                           REGISTERS_0_2_port);
   REGISTERS_reg_0_1_inst : DLH_X1 port map( G => N4592, D => N4533, Q => 
                           REGISTERS_0_1_port);
   REGISTERS_reg_0_0_inst : DLH_X1 port map( G => N4592, D => N4531, Q => 
                           REGISTERS_0_0_port);
   REGISTERS_reg_1_31_inst : DLH_X1 port map( G => N4528, D => N4593, Q => 
                           REGISTERS_1_31_port);
   REGISTERS_reg_1_30_inst : DLH_X1 port map( G => N4528, D => N4591, Q => 
                           REGISTERS_1_30_port);
   REGISTERS_reg_1_29_inst : DLH_X1 port map( G => N4528, D => N4589, Q => 
                           REGISTERS_1_29_port);
   REGISTERS_reg_1_28_inst : DLH_X1 port map( G => N4528, D => N4587, Q => 
                           REGISTERS_1_28_port);
   REGISTERS_reg_1_27_inst : DLH_X1 port map( G => N4528, D => N4585, Q => 
                           REGISTERS_1_27_port);
   REGISTERS_reg_1_26_inst : DLH_X1 port map( G => N4528, D => N4583, Q => 
                           REGISTERS_1_26_port);
   REGISTERS_reg_1_25_inst : DLH_X1 port map( G => N4528, D => N4581, Q => 
                           REGISTERS_1_25_port);
   REGISTERS_reg_1_24_inst : DLH_X1 port map( G => N4528, D => N4579, Q => 
                           REGISTERS_1_24_port);
   REGISTERS_reg_1_23_inst : DLH_X1 port map( G => N4528, D => N4577, Q => 
                           REGISTERS_1_23_port);
   REGISTERS_reg_1_22_inst : DLH_X1 port map( G => N4528, D => N4575, Q => 
                           REGISTERS_1_22_port);
   REGISTERS_reg_1_21_inst : DLH_X1 port map( G => N4528, D => N4573, Q => 
                           REGISTERS_1_21_port);
   REGISTERS_reg_1_20_inst : DLH_X1 port map( G => N4528, D => N4571, Q => 
                           REGISTERS_1_20_port);
   REGISTERS_reg_1_19_inst : DLH_X1 port map( G => N4528, D => N4569, Q => 
                           REGISTERS_1_19_port);
   REGISTERS_reg_1_18_inst : DLH_X1 port map( G => N4528, D => N4567, Q => 
                           REGISTERS_1_18_port);
   REGISTERS_reg_1_17_inst : DLH_X1 port map( G => N4528, D => N4565, Q => 
                           REGISTERS_1_17_port);
   REGISTERS_reg_1_16_inst : DLH_X1 port map( G => N4528, D => N4563, Q => 
                           REGISTERS_1_16_port);
   REGISTERS_reg_1_15_inst : DLH_X1 port map( G => N4528, D => N4561, Q => 
                           REGISTERS_1_15_port);
   REGISTERS_reg_1_14_inst : DLH_X1 port map( G => N4528, D => N4559, Q => 
                           REGISTERS_1_14_port);
   REGISTERS_reg_1_13_inst : DLH_X1 port map( G => N4528, D => N4557, Q => 
                           REGISTERS_1_13_port);
   REGISTERS_reg_1_12_inst : DLH_X1 port map( G => N4528, D => N4555, Q => 
                           REGISTERS_1_12_port);
   REGISTERS_reg_1_11_inst : DLH_X1 port map( G => N4528, D => N4553, Q => 
                           REGISTERS_1_11_port);
   REGISTERS_reg_1_10_inst : DLH_X1 port map( G => N4528, D => N4551, Q => 
                           REGISTERS_1_10_port);
   REGISTERS_reg_1_9_inst : DLH_X1 port map( G => N4528, D => N4549, Q => 
                           REGISTERS_1_9_port);
   REGISTERS_reg_1_8_inst : DLH_X1 port map( G => N4528, D => N4547, Q => 
                           REGISTERS_1_8_port);
   REGISTERS_reg_1_7_inst : DLH_X1 port map( G => N4528, D => N4545, Q => 
                           REGISTERS_1_7_port);
   REGISTERS_reg_1_6_inst : DLH_X1 port map( G => N4528, D => N4543, Q => 
                           REGISTERS_1_6_port);
   REGISTERS_reg_1_5_inst : DLH_X1 port map( G => N4528, D => N4541, Q => 
                           REGISTERS_1_5_port);
   REGISTERS_reg_1_4_inst : DLH_X1 port map( G => N4528, D => N4539, Q => 
                           REGISTERS_1_4_port);
   REGISTERS_reg_1_3_inst : DLH_X1 port map( G => N4528, D => N4537, Q => 
                           REGISTERS_1_3_port);
   REGISTERS_reg_1_2_inst : DLH_X1 port map( G => N4528, D => N4535, Q => 
                           REGISTERS_1_2_port);
   REGISTERS_reg_1_1_inst : DLH_X1 port map( G => N4528, D => N4533, Q => 
                           REGISTERS_1_1_port);
   REGISTERS_reg_1_0_inst : DLH_X1 port map( G => N4528, D => N4531, Q => 
                           REGISTERS_1_0_port);
   REGISTERS_reg_2_31_inst : DLH_X1 port map( G => N4464, D => N4593, Q => 
                           REGISTERS_2_31_port);
   REGISTERS_reg_2_30_inst : DLH_X1 port map( G => N4464, D => N4591, Q => 
                           REGISTERS_2_30_port);
   REGISTERS_reg_2_29_inst : DLH_X1 port map( G => N4464, D => N4589, Q => 
                           REGISTERS_2_29_port);
   REGISTERS_reg_2_28_inst : DLH_X1 port map( G => N4464, D => N4587, Q => 
                           REGISTERS_2_28_port);
   REGISTERS_reg_2_27_inst : DLH_X1 port map( G => N4464, D => N4585, Q => 
                           REGISTERS_2_27_port);
   REGISTERS_reg_2_26_inst : DLH_X1 port map( G => N4464, D => N4583, Q => 
                           REGISTERS_2_26_port);
   REGISTERS_reg_2_25_inst : DLH_X1 port map( G => N4464, D => N4581, Q => 
                           REGISTERS_2_25_port);
   REGISTERS_reg_2_24_inst : DLH_X1 port map( G => N4464, D => N4579, Q => 
                           REGISTERS_2_24_port);
   REGISTERS_reg_2_23_inst : DLH_X1 port map( G => N4464, D => N4577, Q => 
                           REGISTERS_2_23_port);
   REGISTERS_reg_2_22_inst : DLH_X1 port map( G => N4464, D => N4575, Q => 
                           REGISTERS_2_22_port);
   REGISTERS_reg_2_21_inst : DLH_X1 port map( G => N4464, D => N4573, Q => 
                           REGISTERS_2_21_port);
   REGISTERS_reg_2_20_inst : DLH_X1 port map( G => N4464, D => N4571, Q => 
                           REGISTERS_2_20_port);
   REGISTERS_reg_2_19_inst : DLH_X1 port map( G => N4464, D => N4569, Q => 
                           REGISTERS_2_19_port);
   REGISTERS_reg_2_18_inst : DLH_X1 port map( G => N4464, D => N4567, Q => 
                           REGISTERS_2_18_port);
   REGISTERS_reg_2_17_inst : DLH_X1 port map( G => N4464, D => N4565, Q => 
                           REGISTERS_2_17_port);
   REGISTERS_reg_2_16_inst : DLH_X1 port map( G => N4464, D => N4563, Q => 
                           REGISTERS_2_16_port);
   REGISTERS_reg_2_15_inst : DLH_X1 port map( G => N4464, D => N4561, Q => 
                           REGISTERS_2_15_port);
   REGISTERS_reg_2_14_inst : DLH_X1 port map( G => N4464, D => N4559, Q => 
                           REGISTERS_2_14_port);
   REGISTERS_reg_2_13_inst : DLH_X1 port map( G => N4464, D => N4557, Q => 
                           REGISTERS_2_13_port);
   REGISTERS_reg_2_12_inst : DLH_X1 port map( G => N4464, D => N4555, Q => 
                           REGISTERS_2_12_port);
   REGISTERS_reg_2_11_inst : DLH_X1 port map( G => N4464, D => N4553, Q => 
                           REGISTERS_2_11_port);
   REGISTERS_reg_2_10_inst : DLH_X1 port map( G => N4464, D => N4551, Q => 
                           REGISTERS_2_10_port);
   REGISTERS_reg_2_9_inst : DLH_X1 port map( G => N4464, D => N4549, Q => 
                           REGISTERS_2_9_port);
   REGISTERS_reg_2_8_inst : DLH_X1 port map( G => N4464, D => N4547, Q => 
                           REGISTERS_2_8_port);
   REGISTERS_reg_2_7_inst : DLH_X1 port map( G => N4464, D => N4545, Q => 
                           REGISTERS_2_7_port);
   REGISTERS_reg_2_6_inst : DLH_X1 port map( G => N4464, D => N4543, Q => 
                           REGISTERS_2_6_port);
   REGISTERS_reg_2_5_inst : DLH_X1 port map( G => N4464, D => N4541, Q => 
                           REGISTERS_2_5_port);
   REGISTERS_reg_2_4_inst : DLH_X1 port map( G => N4464, D => N4539, Q => 
                           REGISTERS_2_4_port);
   REGISTERS_reg_2_3_inst : DLH_X1 port map( G => N4464, D => N4537, Q => 
                           REGISTERS_2_3_port);
   REGISTERS_reg_2_2_inst : DLH_X1 port map( G => N4464, D => N4535, Q => 
                           REGISTERS_2_2_port);
   REGISTERS_reg_2_1_inst : DLH_X1 port map( G => N4464, D => N4533, Q => 
                           REGISTERS_2_1_port);
   REGISTERS_reg_2_0_inst : DLH_X1 port map( G => N4464, D => N4531, Q => 
                           REGISTERS_2_0_port);
   REGISTERS_reg_3_31_inst : DLH_X1 port map( G => N4400, D => N4593, Q => 
                           REGISTERS_3_31_port);
   REGISTERS_reg_3_30_inst : DLH_X1 port map( G => N4400, D => N4591, Q => 
                           REGISTERS_3_30_port);
   REGISTERS_reg_3_29_inst : DLH_X1 port map( G => N4400, D => N4589, Q => 
                           REGISTERS_3_29_port);
   REGISTERS_reg_3_28_inst : DLH_X1 port map( G => N4400, D => N4587, Q => 
                           REGISTERS_3_28_port);
   REGISTERS_reg_3_27_inst : DLH_X1 port map( G => N4400, D => N4585, Q => 
                           REGISTERS_3_27_port);
   REGISTERS_reg_3_26_inst : DLH_X1 port map( G => N4400, D => N4583, Q => 
                           REGISTERS_3_26_port);
   REGISTERS_reg_3_25_inst : DLH_X1 port map( G => N4400, D => N4581, Q => 
                           REGISTERS_3_25_port);
   REGISTERS_reg_3_24_inst : DLH_X1 port map( G => N4400, D => N4579, Q => 
                           REGISTERS_3_24_port);
   REGISTERS_reg_3_23_inst : DLH_X1 port map( G => N4400, D => N4577, Q => 
                           REGISTERS_3_23_port);
   REGISTERS_reg_3_22_inst : DLH_X1 port map( G => N4400, D => N4575, Q => 
                           REGISTERS_3_22_port);
   REGISTERS_reg_3_21_inst : DLH_X1 port map( G => N4400, D => N4573, Q => 
                           REGISTERS_3_21_port);
   REGISTERS_reg_3_20_inst : DLH_X1 port map( G => N4400, D => N4571, Q => 
                           REGISTERS_3_20_port);
   REGISTERS_reg_3_19_inst : DLH_X1 port map( G => N4400, D => N4569, Q => 
                           REGISTERS_3_19_port);
   REGISTERS_reg_3_18_inst : DLH_X1 port map( G => N4400, D => N4567, Q => 
                           REGISTERS_3_18_port);
   REGISTERS_reg_3_17_inst : DLH_X1 port map( G => N4400, D => N4565, Q => 
                           REGISTERS_3_17_port);
   REGISTERS_reg_3_16_inst : DLH_X1 port map( G => N4400, D => N4563, Q => 
                           REGISTERS_3_16_port);
   REGISTERS_reg_3_15_inst : DLH_X1 port map( G => N4400, D => N4561, Q => 
                           REGISTERS_3_15_port);
   REGISTERS_reg_3_14_inst : DLH_X1 port map( G => N4400, D => N4559, Q => 
                           REGISTERS_3_14_port);
   REGISTERS_reg_3_13_inst : DLH_X1 port map( G => N4400, D => N4557, Q => 
                           REGISTERS_3_13_port);
   REGISTERS_reg_3_12_inst : DLH_X1 port map( G => N4400, D => N4555, Q => 
                           REGISTERS_3_12_port);
   REGISTERS_reg_3_11_inst : DLH_X1 port map( G => N4400, D => N4553, Q => 
                           REGISTERS_3_11_port);
   REGISTERS_reg_3_10_inst : DLH_X1 port map( G => N4400, D => N4551, Q => 
                           REGISTERS_3_10_port);
   REGISTERS_reg_3_9_inst : DLH_X1 port map( G => N4400, D => N4549, Q => 
                           REGISTERS_3_9_port);
   REGISTERS_reg_3_8_inst : DLH_X1 port map( G => N4400, D => N4547, Q => 
                           REGISTERS_3_8_port);
   REGISTERS_reg_3_7_inst : DLH_X1 port map( G => N4400, D => N4545, Q => 
                           REGISTERS_3_7_port);
   REGISTERS_reg_3_6_inst : DLH_X1 port map( G => N4400, D => N4543, Q => 
                           REGISTERS_3_6_port);
   REGISTERS_reg_3_5_inst : DLH_X1 port map( G => N4400, D => N4541, Q => 
                           REGISTERS_3_5_port);
   REGISTERS_reg_3_4_inst : DLH_X1 port map( G => N4400, D => N4539, Q => 
                           REGISTERS_3_4_port);
   REGISTERS_reg_3_3_inst : DLH_X1 port map( G => N4400, D => N4537, Q => 
                           REGISTERS_3_3_port);
   REGISTERS_reg_3_2_inst : DLH_X1 port map( G => N4400, D => N4535, Q => 
                           REGISTERS_3_2_port);
   REGISTERS_reg_3_1_inst : DLH_X1 port map( G => N4400, D => N4533, Q => 
                           REGISTERS_3_1_port);
   REGISTERS_reg_3_0_inst : DLH_X1 port map( G => N4400, D => N4531, Q => 
                           REGISTERS_3_0_port);
   REGISTERS_reg_4_31_inst : DLH_X1 port map( G => N4336, D => N4593, Q => 
                           REGISTERS_4_31_port);
   REGISTERS_reg_4_30_inst : DLH_X1 port map( G => N4336, D => N4591, Q => 
                           REGISTERS_4_30_port);
   REGISTERS_reg_4_29_inst : DLH_X1 port map( G => N4336, D => N4589, Q => 
                           REGISTERS_4_29_port);
   REGISTERS_reg_4_28_inst : DLH_X1 port map( G => N4336, D => N4587, Q => 
                           REGISTERS_4_28_port);
   REGISTERS_reg_4_27_inst : DLH_X1 port map( G => N4336, D => N4585, Q => 
                           REGISTERS_4_27_port);
   REGISTERS_reg_4_26_inst : DLH_X1 port map( G => N4336, D => N4583, Q => 
                           REGISTERS_4_26_port);
   REGISTERS_reg_4_25_inst : DLH_X1 port map( G => N4336, D => N4581, Q => 
                           REGISTERS_4_25_port);
   REGISTERS_reg_4_24_inst : DLH_X1 port map( G => N4336, D => N4579, Q => 
                           REGISTERS_4_24_port);
   REGISTERS_reg_4_23_inst : DLH_X1 port map( G => N4336, D => N4577, Q => 
                           REGISTERS_4_23_port);
   REGISTERS_reg_4_22_inst : DLH_X1 port map( G => N4336, D => N4575, Q => 
                           REGISTERS_4_22_port);
   REGISTERS_reg_4_21_inst : DLH_X1 port map( G => N4336, D => N4573, Q => 
                           REGISTERS_4_21_port);
   REGISTERS_reg_4_20_inst : DLH_X1 port map( G => N4336, D => N4571, Q => 
                           REGISTERS_4_20_port);
   REGISTERS_reg_4_19_inst : DLH_X1 port map( G => N4336, D => N4569, Q => 
                           REGISTERS_4_19_port);
   REGISTERS_reg_4_18_inst : DLH_X1 port map( G => N4336, D => N4567, Q => 
                           REGISTERS_4_18_port);
   REGISTERS_reg_4_17_inst : DLH_X1 port map( G => N4336, D => N4565, Q => 
                           REGISTERS_4_17_port);
   REGISTERS_reg_4_16_inst : DLH_X1 port map( G => N4336, D => N4563, Q => 
                           REGISTERS_4_16_port);
   REGISTERS_reg_4_15_inst : DLH_X1 port map( G => N4336, D => N4561, Q => 
                           REGISTERS_4_15_port);
   REGISTERS_reg_4_14_inst : DLH_X1 port map( G => N4336, D => N4559, Q => 
                           REGISTERS_4_14_port);
   REGISTERS_reg_4_13_inst : DLH_X1 port map( G => N4336, D => N4557, Q => 
                           REGISTERS_4_13_port);
   REGISTERS_reg_4_12_inst : DLH_X1 port map( G => N4336, D => N4555, Q => 
                           REGISTERS_4_12_port);
   REGISTERS_reg_4_11_inst : DLH_X1 port map( G => N4336, D => N4553, Q => 
                           REGISTERS_4_11_port);
   REGISTERS_reg_4_10_inst : DLH_X1 port map( G => N4336, D => N4551, Q => 
                           REGISTERS_4_10_port);
   REGISTERS_reg_4_9_inst : DLH_X1 port map( G => N4336, D => N4549, Q => 
                           REGISTERS_4_9_port);
   REGISTERS_reg_4_8_inst : DLH_X1 port map( G => N4336, D => N4547, Q => 
                           REGISTERS_4_8_port);
   REGISTERS_reg_4_7_inst : DLH_X1 port map( G => N4336, D => N4545, Q => 
                           REGISTERS_4_7_port);
   REGISTERS_reg_4_6_inst : DLH_X1 port map( G => N4336, D => N4543, Q => 
                           REGISTERS_4_6_port);
   REGISTERS_reg_4_5_inst : DLH_X1 port map( G => N4336, D => N4541, Q => 
                           REGISTERS_4_5_port);
   REGISTERS_reg_4_4_inst : DLH_X1 port map( G => N4336, D => N4539, Q => 
                           REGISTERS_4_4_port);
   REGISTERS_reg_4_3_inst : DLH_X1 port map( G => N4336, D => N4537, Q => 
                           REGISTERS_4_3_port);
   REGISTERS_reg_4_2_inst : DLH_X1 port map( G => N4336, D => N4535, Q => 
                           REGISTERS_4_2_port);
   REGISTERS_reg_4_1_inst : DLH_X1 port map( G => N4336, D => N4533, Q => 
                           REGISTERS_4_1_port);
   REGISTERS_reg_4_0_inst : DLH_X1 port map( G => N4336, D => N4531, Q => 
                           REGISTERS_4_0_port);
   REGISTERS_reg_5_31_inst : DLH_X1 port map( G => N4272, D => N4593, Q => 
                           REGISTERS_5_31_port);
   REGISTERS_reg_5_30_inst : DLH_X1 port map( G => N4272, D => N4591, Q => 
                           REGISTERS_5_30_port);
   REGISTERS_reg_5_29_inst : DLH_X1 port map( G => N4272, D => N4589, Q => 
                           REGISTERS_5_29_port);
   REGISTERS_reg_5_28_inst : DLH_X1 port map( G => N4272, D => N4587, Q => 
                           REGISTERS_5_28_port);
   REGISTERS_reg_5_27_inst : DLH_X1 port map( G => N4272, D => N4585, Q => 
                           REGISTERS_5_27_port);
   REGISTERS_reg_5_26_inst : DLH_X1 port map( G => N4272, D => N4583, Q => 
                           REGISTERS_5_26_port);
   REGISTERS_reg_5_25_inst : DLH_X1 port map( G => N4272, D => N4581, Q => 
                           REGISTERS_5_25_port);
   REGISTERS_reg_5_24_inst : DLH_X1 port map( G => N4272, D => N4579, Q => 
                           REGISTERS_5_24_port);
   REGISTERS_reg_5_23_inst : DLH_X1 port map( G => N4272, D => N4577, Q => 
                           REGISTERS_5_23_port);
   REGISTERS_reg_5_22_inst : DLH_X1 port map( G => N4272, D => N4575, Q => 
                           REGISTERS_5_22_port);
   REGISTERS_reg_5_21_inst : DLH_X1 port map( G => N4272, D => N4573, Q => 
                           REGISTERS_5_21_port);
   REGISTERS_reg_5_20_inst : DLH_X1 port map( G => N4272, D => N4571, Q => 
                           REGISTERS_5_20_port);
   REGISTERS_reg_5_19_inst : DLH_X1 port map( G => N4272, D => N4569, Q => 
                           REGISTERS_5_19_port);
   REGISTERS_reg_5_18_inst : DLH_X1 port map( G => N4272, D => N4567, Q => 
                           REGISTERS_5_18_port);
   REGISTERS_reg_5_17_inst : DLH_X1 port map( G => N4272, D => N4565, Q => 
                           REGISTERS_5_17_port);
   REGISTERS_reg_5_16_inst : DLH_X1 port map( G => N4272, D => N4563, Q => 
                           REGISTERS_5_16_port);
   REGISTERS_reg_5_15_inst : DLH_X1 port map( G => N4272, D => N4561, Q => 
                           REGISTERS_5_15_port);
   REGISTERS_reg_5_14_inst : DLH_X1 port map( G => N4272, D => N4559, Q => 
                           REGISTERS_5_14_port);
   REGISTERS_reg_5_13_inst : DLH_X1 port map( G => N4272, D => N4557, Q => 
                           REGISTERS_5_13_port);
   REGISTERS_reg_5_12_inst : DLH_X1 port map( G => N4272, D => N4555, Q => 
                           REGISTERS_5_12_port);
   REGISTERS_reg_5_11_inst : DLH_X1 port map( G => N4272, D => N4553, Q => 
                           REGISTERS_5_11_port);
   REGISTERS_reg_5_10_inst : DLH_X1 port map( G => N4272, D => N4551, Q => 
                           REGISTERS_5_10_port);
   REGISTERS_reg_5_9_inst : DLH_X1 port map( G => N4272, D => N4549, Q => 
                           REGISTERS_5_9_port);
   REGISTERS_reg_5_8_inst : DLH_X1 port map( G => N4272, D => N4547, Q => 
                           REGISTERS_5_8_port);
   REGISTERS_reg_5_7_inst : DLH_X1 port map( G => N4272, D => N4545, Q => 
                           REGISTERS_5_7_port);
   REGISTERS_reg_5_6_inst : DLH_X1 port map( G => N4272, D => N4543, Q => 
                           REGISTERS_5_6_port);
   REGISTERS_reg_5_5_inst : DLH_X1 port map( G => N4272, D => N4541, Q => 
                           REGISTERS_5_5_port);
   REGISTERS_reg_5_4_inst : DLH_X1 port map( G => N4272, D => N4539, Q => 
                           REGISTERS_5_4_port);
   REGISTERS_reg_5_3_inst : DLH_X1 port map( G => N4272, D => N4537, Q => 
                           REGISTERS_5_3_port);
   REGISTERS_reg_5_2_inst : DLH_X1 port map( G => N4272, D => N4535, Q => 
                           REGISTERS_5_2_port);
   REGISTERS_reg_5_1_inst : DLH_X1 port map( G => N4272, D => N4533, Q => 
                           REGISTERS_5_1_port);
   REGISTERS_reg_5_0_inst : DLH_X1 port map( G => N4272, D => N4531, Q => 
                           REGISTERS_5_0_port);
   REGISTERS_reg_6_31_inst : DLH_X1 port map( G => N4208, D => N4593, Q => 
                           REGISTERS_6_31_port);
   REGISTERS_reg_6_30_inst : DLH_X1 port map( G => N4208, D => N4591, Q => 
                           REGISTERS_6_30_port);
   REGISTERS_reg_6_29_inst : DLH_X1 port map( G => N4208, D => N4589, Q => 
                           REGISTERS_6_29_port);
   REGISTERS_reg_6_28_inst : DLH_X1 port map( G => N4208, D => N4587, Q => 
                           REGISTERS_6_28_port);
   REGISTERS_reg_6_27_inst : DLH_X1 port map( G => N4208, D => N4585, Q => 
                           REGISTERS_6_27_port);
   REGISTERS_reg_6_26_inst : DLH_X1 port map( G => N4208, D => N4583, Q => 
                           REGISTERS_6_26_port);
   REGISTERS_reg_6_25_inst : DLH_X1 port map( G => N4208, D => N4581, Q => 
                           REGISTERS_6_25_port);
   REGISTERS_reg_6_24_inst : DLH_X1 port map( G => N4208, D => N4579, Q => 
                           REGISTERS_6_24_port);
   REGISTERS_reg_6_23_inst : DLH_X1 port map( G => N4208, D => N4577, Q => 
                           REGISTERS_6_23_port);
   REGISTERS_reg_6_22_inst : DLH_X1 port map( G => N4208, D => N4575, Q => 
                           REGISTERS_6_22_port);
   REGISTERS_reg_6_21_inst : DLH_X1 port map( G => N4208, D => N4573, Q => 
                           REGISTERS_6_21_port);
   REGISTERS_reg_6_20_inst : DLH_X1 port map( G => N4208, D => N4571, Q => 
                           REGISTERS_6_20_port);
   REGISTERS_reg_6_19_inst : DLH_X1 port map( G => N4208, D => N4569, Q => 
                           REGISTERS_6_19_port);
   REGISTERS_reg_6_18_inst : DLH_X1 port map( G => N4208, D => N4567, Q => 
                           REGISTERS_6_18_port);
   REGISTERS_reg_6_17_inst : DLH_X1 port map( G => N4208, D => N4565, Q => 
                           REGISTERS_6_17_port);
   REGISTERS_reg_6_16_inst : DLH_X1 port map( G => N4208, D => N4563, Q => 
                           REGISTERS_6_16_port);
   REGISTERS_reg_6_15_inst : DLH_X1 port map( G => N4208, D => N4561, Q => 
                           REGISTERS_6_15_port);
   REGISTERS_reg_6_14_inst : DLH_X1 port map( G => N4208, D => N4559, Q => 
                           REGISTERS_6_14_port);
   REGISTERS_reg_6_13_inst : DLH_X1 port map( G => N4208, D => N4557, Q => 
                           REGISTERS_6_13_port);
   REGISTERS_reg_6_12_inst : DLH_X1 port map( G => N4208, D => N4555, Q => 
                           REGISTERS_6_12_port);
   REGISTERS_reg_6_11_inst : DLH_X1 port map( G => N4208, D => N4553, Q => 
                           REGISTERS_6_11_port);
   REGISTERS_reg_6_10_inst : DLH_X1 port map( G => N4208, D => N4551, Q => 
                           REGISTERS_6_10_port);
   REGISTERS_reg_6_9_inst : DLH_X1 port map( G => N4208, D => N4549, Q => 
                           REGISTERS_6_9_port);
   REGISTERS_reg_6_8_inst : DLH_X1 port map( G => N4208, D => N4547, Q => 
                           REGISTERS_6_8_port);
   REGISTERS_reg_6_7_inst : DLH_X1 port map( G => N4208, D => N4545, Q => 
                           REGISTERS_6_7_port);
   REGISTERS_reg_6_6_inst : DLH_X1 port map( G => N4208, D => N4543, Q => 
                           REGISTERS_6_6_port);
   REGISTERS_reg_6_5_inst : DLH_X1 port map( G => N4208, D => N4541, Q => 
                           REGISTERS_6_5_port);
   REGISTERS_reg_6_4_inst : DLH_X1 port map( G => N4208, D => N4539, Q => 
                           REGISTERS_6_4_port);
   REGISTERS_reg_6_3_inst : DLH_X1 port map( G => N4208, D => N4537, Q => 
                           REGISTERS_6_3_port);
   REGISTERS_reg_6_2_inst : DLH_X1 port map( G => N4208, D => N4535, Q => 
                           REGISTERS_6_2_port);
   REGISTERS_reg_6_1_inst : DLH_X1 port map( G => N4208, D => N4533, Q => 
                           REGISTERS_6_1_port);
   REGISTERS_reg_6_0_inst : DLH_X1 port map( G => N4208, D => N4531, Q => 
                           REGISTERS_6_0_port);
   REGISTERS_reg_7_31_inst : DLH_X1 port map( G => N4144, D => N4593, Q => 
                           REGISTERS_7_31_port);
   REGISTERS_reg_7_30_inst : DLH_X1 port map( G => N4144, D => N4591, Q => 
                           REGISTERS_7_30_port);
   REGISTERS_reg_7_29_inst : DLH_X1 port map( G => N4144, D => N4589, Q => 
                           REGISTERS_7_29_port);
   REGISTERS_reg_7_28_inst : DLH_X1 port map( G => N4144, D => N4587, Q => 
                           REGISTERS_7_28_port);
   REGISTERS_reg_7_27_inst : DLH_X1 port map( G => N4144, D => N4585, Q => 
                           REGISTERS_7_27_port);
   REGISTERS_reg_7_26_inst : DLH_X1 port map( G => N4144, D => N4583, Q => 
                           REGISTERS_7_26_port);
   REGISTERS_reg_7_25_inst : DLH_X1 port map( G => N4144, D => N4581, Q => 
                           REGISTERS_7_25_port);
   REGISTERS_reg_7_24_inst : DLH_X1 port map( G => N4144, D => N4579, Q => 
                           REGISTERS_7_24_port);
   REGISTERS_reg_7_23_inst : DLH_X1 port map( G => N4144, D => N4577, Q => 
                           REGISTERS_7_23_port);
   REGISTERS_reg_7_22_inst : DLH_X1 port map( G => N4144, D => N4575, Q => 
                           REGISTERS_7_22_port);
   REGISTERS_reg_7_21_inst : DLH_X1 port map( G => N4144, D => N4573, Q => 
                           REGISTERS_7_21_port);
   REGISTERS_reg_7_20_inst : DLH_X1 port map( G => N4144, D => N4571, Q => 
                           REGISTERS_7_20_port);
   REGISTERS_reg_7_19_inst : DLH_X1 port map( G => N4144, D => N4569, Q => 
                           REGISTERS_7_19_port);
   REGISTERS_reg_7_18_inst : DLH_X1 port map( G => N4144, D => N4567, Q => 
                           REGISTERS_7_18_port);
   REGISTERS_reg_7_17_inst : DLH_X1 port map( G => N4144, D => N4565, Q => 
                           REGISTERS_7_17_port);
   REGISTERS_reg_7_16_inst : DLH_X1 port map( G => N4144, D => N4563, Q => 
                           REGISTERS_7_16_port);
   REGISTERS_reg_7_15_inst : DLH_X1 port map( G => N4144, D => N4561, Q => 
                           REGISTERS_7_15_port);
   REGISTERS_reg_7_14_inst : DLH_X1 port map( G => N4144, D => N4559, Q => 
                           REGISTERS_7_14_port);
   REGISTERS_reg_7_13_inst : DLH_X1 port map( G => N4144, D => N4557, Q => 
                           REGISTERS_7_13_port);
   REGISTERS_reg_7_12_inst : DLH_X1 port map( G => N4144, D => N4555, Q => 
                           REGISTERS_7_12_port);
   REGISTERS_reg_7_11_inst : DLH_X1 port map( G => N4144, D => N4553, Q => 
                           REGISTERS_7_11_port);
   REGISTERS_reg_7_10_inst : DLH_X1 port map( G => N4144, D => N4551, Q => 
                           REGISTERS_7_10_port);
   REGISTERS_reg_7_9_inst : DLH_X1 port map( G => N4144, D => N4549, Q => 
                           REGISTERS_7_9_port);
   REGISTERS_reg_7_8_inst : DLH_X1 port map( G => N4144, D => N4547, Q => 
                           REGISTERS_7_8_port);
   REGISTERS_reg_7_7_inst : DLH_X1 port map( G => N4144, D => N4545, Q => 
                           REGISTERS_7_7_port);
   REGISTERS_reg_7_6_inst : DLH_X1 port map( G => N4144, D => N4543, Q => 
                           REGISTERS_7_6_port);
   REGISTERS_reg_7_5_inst : DLH_X1 port map( G => N4144, D => N4541, Q => 
                           REGISTERS_7_5_port);
   REGISTERS_reg_7_4_inst : DLH_X1 port map( G => N4144, D => N4539, Q => 
                           REGISTERS_7_4_port);
   REGISTERS_reg_7_3_inst : DLH_X1 port map( G => N4144, D => N4537, Q => 
                           REGISTERS_7_3_port);
   REGISTERS_reg_7_2_inst : DLH_X1 port map( G => N4144, D => N4535, Q => 
                           REGISTERS_7_2_port);
   REGISTERS_reg_7_1_inst : DLH_X1 port map( G => N4144, D => N4533, Q => 
                           REGISTERS_7_1_port);
   REGISTERS_reg_7_0_inst : DLH_X1 port map( G => N4144, D => N4531, Q => 
                           REGISTERS_7_0_port);
   REGISTERS_reg_8_31_inst : DLH_X1 port map( G => N4080, D => N4593, Q => 
                           REGISTERS_8_31_port);
   REGISTERS_reg_8_30_inst : DLH_X1 port map( G => N4080, D => N4591, Q => 
                           REGISTERS_8_30_port);
   REGISTERS_reg_8_29_inst : DLH_X1 port map( G => N4080, D => N4589, Q => 
                           REGISTERS_8_29_port);
   REGISTERS_reg_8_28_inst : DLH_X1 port map( G => N4080, D => N4587, Q => 
                           REGISTERS_8_28_port);
   REGISTERS_reg_8_27_inst : DLH_X1 port map( G => N4080, D => N4585, Q => 
                           REGISTERS_8_27_port);
   REGISTERS_reg_8_26_inst : DLH_X1 port map( G => N4080, D => N4583, Q => 
                           REGISTERS_8_26_port);
   REGISTERS_reg_8_25_inst : DLH_X1 port map( G => N4080, D => N4581, Q => 
                           REGISTERS_8_25_port);
   REGISTERS_reg_8_24_inst : DLH_X1 port map( G => N4080, D => N4579, Q => 
                           REGISTERS_8_24_port);
   REGISTERS_reg_8_23_inst : DLH_X1 port map( G => N4080, D => N4577, Q => 
                           REGISTERS_8_23_port);
   REGISTERS_reg_8_22_inst : DLH_X1 port map( G => N4080, D => N4575, Q => 
                           REGISTERS_8_22_port);
   REGISTERS_reg_8_21_inst : DLH_X1 port map( G => N4080, D => N4573, Q => 
                           REGISTERS_8_21_port);
   REGISTERS_reg_8_20_inst : DLH_X1 port map( G => N4080, D => N4571, Q => 
                           REGISTERS_8_20_port);
   REGISTERS_reg_8_19_inst : DLH_X1 port map( G => N4080, D => N4569, Q => 
                           REGISTERS_8_19_port);
   REGISTERS_reg_8_18_inst : DLH_X1 port map( G => N4080, D => N4567, Q => 
                           REGISTERS_8_18_port);
   REGISTERS_reg_8_17_inst : DLH_X1 port map( G => N4080, D => N4565, Q => 
                           REGISTERS_8_17_port);
   REGISTERS_reg_8_16_inst : DLH_X1 port map( G => N4080, D => N4563, Q => 
                           REGISTERS_8_16_port);
   REGISTERS_reg_8_15_inst : DLH_X1 port map( G => N4080, D => N4561, Q => 
                           REGISTERS_8_15_port);
   REGISTERS_reg_8_14_inst : DLH_X1 port map( G => N4080, D => N4559, Q => 
                           REGISTERS_8_14_port);
   REGISTERS_reg_8_13_inst : DLH_X1 port map( G => N4080, D => N4557, Q => 
                           REGISTERS_8_13_port);
   REGISTERS_reg_8_12_inst : DLH_X1 port map( G => N4080, D => N4555, Q => 
                           REGISTERS_8_12_port);
   REGISTERS_reg_8_11_inst : DLH_X1 port map( G => N4080, D => N4553, Q => 
                           REGISTERS_8_11_port);
   REGISTERS_reg_8_10_inst : DLH_X1 port map( G => N4080, D => N4551, Q => 
                           REGISTERS_8_10_port);
   REGISTERS_reg_8_9_inst : DLH_X1 port map( G => N4080, D => N4549, Q => 
                           REGISTERS_8_9_port);
   REGISTERS_reg_8_8_inst : DLH_X1 port map( G => N4080, D => N4547, Q => 
                           REGISTERS_8_8_port);
   REGISTERS_reg_8_7_inst : DLH_X1 port map( G => N4080, D => N4545, Q => 
                           REGISTERS_8_7_port);
   REGISTERS_reg_8_6_inst : DLH_X1 port map( G => N4080, D => N4543, Q => 
                           REGISTERS_8_6_port);
   REGISTERS_reg_8_5_inst : DLH_X1 port map( G => N4080, D => N4541, Q => 
                           REGISTERS_8_5_port);
   REGISTERS_reg_8_4_inst : DLH_X1 port map( G => N4080, D => N4539, Q => 
                           REGISTERS_8_4_port);
   REGISTERS_reg_8_3_inst : DLH_X1 port map( G => N4080, D => N4537, Q => 
                           REGISTERS_8_3_port);
   REGISTERS_reg_8_2_inst : DLH_X1 port map( G => N4080, D => N4535, Q => 
                           REGISTERS_8_2_port);
   REGISTERS_reg_8_1_inst : DLH_X1 port map( G => N4080, D => N4533, Q => 
                           REGISTERS_8_1_port);
   REGISTERS_reg_8_0_inst : DLH_X1 port map( G => N4080, D => N4531, Q => 
                           REGISTERS_8_0_port);
   REGISTERS_reg_9_31_inst : DLH_X1 port map( G => N4016, D => N4593, Q => 
                           REGISTERS_9_31_port);
   REGISTERS_reg_9_30_inst : DLH_X1 port map( G => N4016, D => N4591, Q => 
                           REGISTERS_9_30_port);
   REGISTERS_reg_9_29_inst : DLH_X1 port map( G => N4016, D => N4589, Q => 
                           REGISTERS_9_29_port);
   REGISTERS_reg_9_28_inst : DLH_X1 port map( G => N4016, D => N4587, Q => 
                           REGISTERS_9_28_port);
   REGISTERS_reg_9_27_inst : DLH_X1 port map( G => N4016, D => N4585, Q => 
                           REGISTERS_9_27_port);
   REGISTERS_reg_9_26_inst : DLH_X1 port map( G => N4016, D => N4583, Q => 
                           REGISTERS_9_26_port);
   REGISTERS_reg_9_25_inst : DLH_X1 port map( G => N4016, D => N4581, Q => 
                           REGISTERS_9_25_port);
   REGISTERS_reg_9_24_inst : DLH_X1 port map( G => N4016, D => N4579, Q => 
                           REGISTERS_9_24_port);
   REGISTERS_reg_9_23_inst : DLH_X1 port map( G => N4016, D => N4577, Q => 
                           REGISTERS_9_23_port);
   REGISTERS_reg_9_22_inst : DLH_X1 port map( G => N4016, D => N4575, Q => 
                           REGISTERS_9_22_port);
   REGISTERS_reg_9_21_inst : DLH_X1 port map( G => N4016, D => N4573, Q => 
                           REGISTERS_9_21_port);
   REGISTERS_reg_9_20_inst : DLH_X1 port map( G => N4016, D => N4571, Q => 
                           REGISTERS_9_20_port);
   REGISTERS_reg_9_19_inst : DLH_X1 port map( G => N4016, D => N4569, Q => 
                           REGISTERS_9_19_port);
   REGISTERS_reg_9_18_inst : DLH_X1 port map( G => N4016, D => N4567, Q => 
                           REGISTERS_9_18_port);
   REGISTERS_reg_9_17_inst : DLH_X1 port map( G => N4016, D => N4565, Q => 
                           REGISTERS_9_17_port);
   REGISTERS_reg_9_16_inst : DLH_X1 port map( G => N4016, D => N4563, Q => 
                           REGISTERS_9_16_port);
   REGISTERS_reg_9_15_inst : DLH_X1 port map( G => N4016, D => N4561, Q => 
                           REGISTERS_9_15_port);
   REGISTERS_reg_9_14_inst : DLH_X1 port map( G => N4016, D => N4559, Q => 
                           REGISTERS_9_14_port);
   REGISTERS_reg_9_13_inst : DLH_X1 port map( G => N4016, D => N4557, Q => 
                           REGISTERS_9_13_port);
   REGISTERS_reg_9_12_inst : DLH_X1 port map( G => N4016, D => N4555, Q => 
                           REGISTERS_9_12_port);
   REGISTERS_reg_9_11_inst : DLH_X1 port map( G => N4016, D => N4553, Q => 
                           REGISTERS_9_11_port);
   REGISTERS_reg_9_10_inst : DLH_X1 port map( G => N4016, D => N4551, Q => 
                           REGISTERS_9_10_port);
   REGISTERS_reg_9_9_inst : DLH_X1 port map( G => N4016, D => N4549, Q => 
                           REGISTERS_9_9_port);
   REGISTERS_reg_9_8_inst : DLH_X1 port map( G => N4016, D => N4547, Q => 
                           REGISTERS_9_8_port);
   REGISTERS_reg_9_7_inst : DLH_X1 port map( G => N4016, D => N4545, Q => 
                           REGISTERS_9_7_port);
   REGISTERS_reg_9_6_inst : DLH_X1 port map( G => N4016, D => N4543, Q => 
                           REGISTERS_9_6_port);
   REGISTERS_reg_9_5_inst : DLH_X1 port map( G => N4016, D => N4541, Q => 
                           REGISTERS_9_5_port);
   REGISTERS_reg_9_4_inst : DLH_X1 port map( G => N4016, D => N4539, Q => 
                           REGISTERS_9_4_port);
   REGISTERS_reg_9_3_inst : DLH_X1 port map( G => N4016, D => N4537, Q => 
                           REGISTERS_9_3_port);
   REGISTERS_reg_9_2_inst : DLH_X1 port map( G => N4016, D => N4535, Q => 
                           REGISTERS_9_2_port);
   REGISTERS_reg_9_1_inst : DLH_X1 port map( G => N4016, D => N4533, Q => 
                           REGISTERS_9_1_port);
   REGISTERS_reg_9_0_inst : DLH_X1 port map( G => N4016, D => N4531, Q => 
                           REGISTERS_9_0_port);
   REGISTERS_reg_10_31_inst : DLH_X1 port map( G => N3952, D => N4593, Q => 
                           REGISTERS_10_31_port);
   REGISTERS_reg_10_30_inst : DLH_X1 port map( G => N3952, D => N4591, Q => 
                           REGISTERS_10_30_port);
   REGISTERS_reg_10_29_inst : DLH_X1 port map( G => N3952, D => N4589, Q => 
                           REGISTERS_10_29_port);
   REGISTERS_reg_10_28_inst : DLH_X1 port map( G => N3952, D => N4587, Q => 
                           REGISTERS_10_28_port);
   REGISTERS_reg_10_27_inst : DLH_X1 port map( G => N3952, D => N4585, Q => 
                           REGISTERS_10_27_port);
   REGISTERS_reg_10_26_inst : DLH_X1 port map( G => N3952, D => N4583, Q => 
                           REGISTERS_10_26_port);
   REGISTERS_reg_10_25_inst : DLH_X1 port map( G => N3952, D => N4581, Q => 
                           REGISTERS_10_25_port);
   REGISTERS_reg_10_24_inst : DLH_X1 port map( G => N3952, D => N4579, Q => 
                           REGISTERS_10_24_port);
   REGISTERS_reg_10_23_inst : DLH_X1 port map( G => N3952, D => N4577, Q => 
                           REGISTERS_10_23_port);
   REGISTERS_reg_10_22_inst : DLH_X1 port map( G => N3952, D => N4575, Q => 
                           REGISTERS_10_22_port);
   REGISTERS_reg_10_21_inst : DLH_X1 port map( G => N3952, D => N4573, Q => 
                           REGISTERS_10_21_port);
   REGISTERS_reg_10_20_inst : DLH_X1 port map( G => N3952, D => N4571, Q => 
                           REGISTERS_10_20_port);
   REGISTERS_reg_10_19_inst : DLH_X1 port map( G => N3952, D => N4569, Q => 
                           REGISTERS_10_19_port);
   REGISTERS_reg_10_18_inst : DLH_X1 port map( G => N3952, D => N4567, Q => 
                           REGISTERS_10_18_port);
   REGISTERS_reg_10_17_inst : DLH_X1 port map( G => N3952, D => N4565, Q => 
                           REGISTERS_10_17_port);
   REGISTERS_reg_10_16_inst : DLH_X1 port map( G => N3952, D => N4563, Q => 
                           REGISTERS_10_16_port);
   REGISTERS_reg_10_15_inst : DLH_X1 port map( G => N3952, D => N4561, Q => 
                           REGISTERS_10_15_port);
   REGISTERS_reg_10_14_inst : DLH_X1 port map( G => N3952, D => N4559, Q => 
                           REGISTERS_10_14_port);
   REGISTERS_reg_10_13_inst : DLH_X1 port map( G => N3952, D => N4557, Q => 
                           REGISTERS_10_13_port);
   REGISTERS_reg_10_12_inst : DLH_X1 port map( G => N3952, D => N4555, Q => 
                           REGISTERS_10_12_port);
   REGISTERS_reg_10_11_inst : DLH_X1 port map( G => N3952, D => N4553, Q => 
                           REGISTERS_10_11_port);
   REGISTERS_reg_10_10_inst : DLH_X1 port map( G => N3952, D => N4551, Q => 
                           REGISTERS_10_10_port);
   REGISTERS_reg_10_9_inst : DLH_X1 port map( G => N3952, D => N4549, Q => 
                           REGISTERS_10_9_port);
   REGISTERS_reg_10_8_inst : DLH_X1 port map( G => N3952, D => N4547, Q => 
                           REGISTERS_10_8_port);
   REGISTERS_reg_10_7_inst : DLH_X1 port map( G => N3952, D => N4545, Q => 
                           REGISTERS_10_7_port);
   REGISTERS_reg_10_6_inst : DLH_X1 port map( G => N3952, D => N4543, Q => 
                           REGISTERS_10_6_port);
   REGISTERS_reg_10_5_inst : DLH_X1 port map( G => N3952, D => N4541, Q => 
                           REGISTERS_10_5_port);
   REGISTERS_reg_10_4_inst : DLH_X1 port map( G => N3952, D => N4539, Q => 
                           REGISTERS_10_4_port);
   REGISTERS_reg_10_3_inst : DLH_X1 port map( G => N3952, D => N4537, Q => 
                           REGISTERS_10_3_port);
   REGISTERS_reg_10_2_inst : DLH_X1 port map( G => N3952, D => N4535, Q => 
                           REGISTERS_10_2_port);
   REGISTERS_reg_10_1_inst : DLH_X1 port map( G => N3952, D => N4533, Q => 
                           REGISTERS_10_1_port);
   REGISTERS_reg_10_0_inst : DLH_X1 port map( G => N3952, D => N4531, Q => 
                           REGISTERS_10_0_port);
   REGISTERS_reg_11_31_inst : DLH_X1 port map( G => N3888, D => N4593, Q => 
                           REGISTERS_11_31_port);
   REGISTERS_reg_11_30_inst : DLH_X1 port map( G => N3888, D => N4591, Q => 
                           REGISTERS_11_30_port);
   REGISTERS_reg_11_29_inst : DLH_X1 port map( G => N3888, D => N4589, Q => 
                           REGISTERS_11_29_port);
   REGISTERS_reg_11_28_inst : DLH_X1 port map( G => N3888, D => N4587, Q => 
                           REGISTERS_11_28_port);
   REGISTERS_reg_11_27_inst : DLH_X1 port map( G => N3888, D => N4585, Q => 
                           REGISTERS_11_27_port);
   REGISTERS_reg_11_26_inst : DLH_X1 port map( G => N3888, D => N4583, Q => 
                           REGISTERS_11_26_port);
   REGISTERS_reg_11_25_inst : DLH_X1 port map( G => N3888, D => N4581, Q => 
                           REGISTERS_11_25_port);
   REGISTERS_reg_11_24_inst : DLH_X1 port map( G => N3888, D => N4579, Q => 
                           REGISTERS_11_24_port);
   REGISTERS_reg_11_23_inst : DLH_X1 port map( G => N3888, D => N4577, Q => 
                           REGISTERS_11_23_port);
   REGISTERS_reg_11_22_inst : DLH_X1 port map( G => N3888, D => N4575, Q => 
                           REGISTERS_11_22_port);
   REGISTERS_reg_11_21_inst : DLH_X1 port map( G => N3888, D => N4573, Q => 
                           REGISTERS_11_21_port);
   REGISTERS_reg_11_20_inst : DLH_X1 port map( G => N3888, D => N4571, Q => 
                           REGISTERS_11_20_port);
   REGISTERS_reg_11_19_inst : DLH_X1 port map( G => N3888, D => N4569, Q => 
                           REGISTERS_11_19_port);
   REGISTERS_reg_11_18_inst : DLH_X1 port map( G => N3888, D => N4567, Q => 
                           REGISTERS_11_18_port);
   REGISTERS_reg_11_17_inst : DLH_X1 port map( G => N3888, D => N4565, Q => 
                           REGISTERS_11_17_port);
   REGISTERS_reg_11_16_inst : DLH_X1 port map( G => N3888, D => N4563, Q => 
                           REGISTERS_11_16_port);
   REGISTERS_reg_11_15_inst : DLH_X1 port map( G => N3888, D => N4561, Q => 
                           REGISTERS_11_15_port);
   REGISTERS_reg_11_14_inst : DLH_X1 port map( G => N3888, D => N4559, Q => 
                           REGISTERS_11_14_port);
   REGISTERS_reg_11_13_inst : DLH_X1 port map( G => N3888, D => N4557, Q => 
                           REGISTERS_11_13_port);
   REGISTERS_reg_11_12_inst : DLH_X1 port map( G => N3888, D => N4555, Q => 
                           REGISTERS_11_12_port);
   REGISTERS_reg_11_11_inst : DLH_X1 port map( G => N3888, D => N4553, Q => 
                           REGISTERS_11_11_port);
   REGISTERS_reg_11_10_inst : DLH_X1 port map( G => N3888, D => N4551, Q => 
                           REGISTERS_11_10_port);
   REGISTERS_reg_11_9_inst : DLH_X1 port map( G => N3888, D => N4549, Q => 
                           REGISTERS_11_9_port);
   REGISTERS_reg_11_8_inst : DLH_X1 port map( G => N3888, D => N4547, Q => 
                           REGISTERS_11_8_port);
   REGISTERS_reg_11_7_inst : DLH_X1 port map( G => N3888, D => N4545, Q => 
                           REGISTERS_11_7_port);
   REGISTERS_reg_11_6_inst : DLH_X1 port map( G => N3888, D => N4543, Q => 
                           REGISTERS_11_6_port);
   REGISTERS_reg_11_5_inst : DLH_X1 port map( G => N3888, D => N4541, Q => 
                           REGISTERS_11_5_port);
   REGISTERS_reg_11_4_inst : DLH_X1 port map( G => N3888, D => N4539, Q => 
                           REGISTERS_11_4_port);
   REGISTERS_reg_11_3_inst : DLH_X1 port map( G => N3888, D => N4537, Q => 
                           REGISTERS_11_3_port);
   REGISTERS_reg_11_2_inst : DLH_X1 port map( G => N3888, D => N4535, Q => 
                           REGISTERS_11_2_port);
   REGISTERS_reg_11_1_inst : DLH_X1 port map( G => N3888, D => N4533, Q => 
                           REGISTERS_11_1_port);
   REGISTERS_reg_11_0_inst : DLH_X1 port map( G => N3888, D => N4531, Q => 
                           REGISTERS_11_0_port);
   REGISTERS_reg_12_31_inst : DLH_X1 port map( G => N3824, D => N4593, Q => 
                           REGISTERS_12_31_port);
   REGISTERS_reg_12_30_inst : DLH_X1 port map( G => N3824, D => N4591, Q => 
                           REGISTERS_12_30_port);
   REGISTERS_reg_12_29_inst : DLH_X1 port map( G => N3824, D => N4589, Q => 
                           REGISTERS_12_29_port);
   REGISTERS_reg_12_28_inst : DLH_X1 port map( G => N3824, D => N4587, Q => 
                           REGISTERS_12_28_port);
   REGISTERS_reg_12_27_inst : DLH_X1 port map( G => N3824, D => N4585, Q => 
                           REGISTERS_12_27_port);
   REGISTERS_reg_12_26_inst : DLH_X1 port map( G => N3824, D => N4583, Q => 
                           REGISTERS_12_26_port);
   REGISTERS_reg_12_25_inst : DLH_X1 port map( G => N3824, D => N4581, Q => 
                           REGISTERS_12_25_port);
   REGISTERS_reg_12_24_inst : DLH_X1 port map( G => N3824, D => N4579, Q => 
                           REGISTERS_12_24_port);
   REGISTERS_reg_12_23_inst : DLH_X1 port map( G => N3824, D => N4577, Q => 
                           REGISTERS_12_23_port);
   REGISTERS_reg_12_22_inst : DLH_X1 port map( G => N3824, D => N4575, Q => 
                           REGISTERS_12_22_port);
   REGISTERS_reg_12_21_inst : DLH_X1 port map( G => N3824, D => N4573, Q => 
                           REGISTERS_12_21_port);
   REGISTERS_reg_12_20_inst : DLH_X1 port map( G => N3824, D => N4571, Q => 
                           REGISTERS_12_20_port);
   REGISTERS_reg_12_19_inst : DLH_X1 port map( G => N3824, D => N4569, Q => 
                           REGISTERS_12_19_port);
   REGISTERS_reg_12_18_inst : DLH_X1 port map( G => N3824, D => N4567, Q => 
                           REGISTERS_12_18_port);
   REGISTERS_reg_12_17_inst : DLH_X1 port map( G => N3824, D => N4565, Q => 
                           REGISTERS_12_17_port);
   REGISTERS_reg_12_16_inst : DLH_X1 port map( G => N3824, D => N4563, Q => 
                           REGISTERS_12_16_port);
   REGISTERS_reg_12_15_inst : DLH_X1 port map( G => N3824, D => N4561, Q => 
                           REGISTERS_12_15_port);
   REGISTERS_reg_12_14_inst : DLH_X1 port map( G => N3824, D => N4559, Q => 
                           REGISTERS_12_14_port);
   REGISTERS_reg_12_13_inst : DLH_X1 port map( G => N3824, D => N4557, Q => 
                           REGISTERS_12_13_port);
   REGISTERS_reg_12_12_inst : DLH_X1 port map( G => N3824, D => N4555, Q => 
                           REGISTERS_12_12_port);
   REGISTERS_reg_12_11_inst : DLH_X1 port map( G => N3824, D => N4553, Q => 
                           REGISTERS_12_11_port);
   REGISTERS_reg_12_10_inst : DLH_X1 port map( G => N3824, D => N4551, Q => 
                           REGISTERS_12_10_port);
   REGISTERS_reg_12_9_inst : DLH_X1 port map( G => N3824, D => N4549, Q => 
                           REGISTERS_12_9_port);
   REGISTERS_reg_12_8_inst : DLH_X1 port map( G => N3824, D => N4547, Q => 
                           REGISTERS_12_8_port);
   REGISTERS_reg_12_7_inst : DLH_X1 port map( G => N3824, D => N4545, Q => 
                           REGISTERS_12_7_port);
   REGISTERS_reg_12_6_inst : DLH_X1 port map( G => N3824, D => N4543, Q => 
                           REGISTERS_12_6_port);
   REGISTERS_reg_12_5_inst : DLH_X1 port map( G => N3824, D => N4541, Q => 
                           REGISTERS_12_5_port);
   REGISTERS_reg_12_4_inst : DLH_X1 port map( G => N3824, D => N4539, Q => 
                           REGISTERS_12_4_port);
   REGISTERS_reg_12_3_inst : DLH_X1 port map( G => N3824, D => N4537, Q => 
                           REGISTERS_12_3_port);
   REGISTERS_reg_12_2_inst : DLH_X1 port map( G => N3824, D => N4535, Q => 
                           REGISTERS_12_2_port);
   REGISTERS_reg_12_1_inst : DLH_X1 port map( G => N3824, D => N4533, Q => 
                           REGISTERS_12_1_port);
   REGISTERS_reg_12_0_inst : DLH_X1 port map( G => N3824, D => N4531, Q => 
                           REGISTERS_12_0_port);
   REGISTERS_reg_13_31_inst : DLH_X1 port map( G => N3760, D => N4593, Q => 
                           REGISTERS_13_31_port);
   REGISTERS_reg_13_30_inst : DLH_X1 port map( G => N3760, D => N4591, Q => 
                           REGISTERS_13_30_port);
   REGISTERS_reg_13_29_inst : DLH_X1 port map( G => N3760, D => N4589, Q => 
                           REGISTERS_13_29_port);
   REGISTERS_reg_13_28_inst : DLH_X1 port map( G => N3760, D => N4587, Q => 
                           REGISTERS_13_28_port);
   REGISTERS_reg_13_27_inst : DLH_X1 port map( G => N3760, D => N4585, Q => 
                           REGISTERS_13_27_port);
   REGISTERS_reg_13_26_inst : DLH_X1 port map( G => N3760, D => N4583, Q => 
                           REGISTERS_13_26_port);
   REGISTERS_reg_13_25_inst : DLH_X1 port map( G => N3760, D => N4581, Q => 
                           REGISTERS_13_25_port);
   REGISTERS_reg_13_24_inst : DLH_X1 port map( G => N3760, D => N4579, Q => 
                           REGISTERS_13_24_port);
   REGISTERS_reg_13_23_inst : DLH_X1 port map( G => N3760, D => N4577, Q => 
                           REGISTERS_13_23_port);
   REGISTERS_reg_13_22_inst : DLH_X1 port map( G => N3760, D => N4575, Q => 
                           REGISTERS_13_22_port);
   REGISTERS_reg_13_21_inst : DLH_X1 port map( G => N3760, D => N4573, Q => 
                           REGISTERS_13_21_port);
   REGISTERS_reg_13_20_inst : DLH_X1 port map( G => N3760, D => N4571, Q => 
                           REGISTERS_13_20_port);
   REGISTERS_reg_13_19_inst : DLH_X1 port map( G => N3760, D => N4569, Q => 
                           REGISTERS_13_19_port);
   REGISTERS_reg_13_18_inst : DLH_X1 port map( G => N3760, D => N4567, Q => 
                           REGISTERS_13_18_port);
   REGISTERS_reg_13_17_inst : DLH_X1 port map( G => N3760, D => N4565, Q => 
                           REGISTERS_13_17_port);
   REGISTERS_reg_13_16_inst : DLH_X1 port map( G => N3760, D => N4563, Q => 
                           REGISTERS_13_16_port);
   REGISTERS_reg_13_15_inst : DLH_X1 port map( G => N3760, D => N4561, Q => 
                           REGISTERS_13_15_port);
   REGISTERS_reg_13_14_inst : DLH_X1 port map( G => N3760, D => N4559, Q => 
                           REGISTERS_13_14_port);
   REGISTERS_reg_13_13_inst : DLH_X1 port map( G => N3760, D => N4557, Q => 
                           REGISTERS_13_13_port);
   REGISTERS_reg_13_12_inst : DLH_X1 port map( G => N3760, D => N4555, Q => 
                           REGISTERS_13_12_port);
   REGISTERS_reg_13_11_inst : DLH_X1 port map( G => N3760, D => N4553, Q => 
                           REGISTERS_13_11_port);
   REGISTERS_reg_13_10_inst : DLH_X1 port map( G => N3760, D => N4551, Q => 
                           REGISTERS_13_10_port);
   REGISTERS_reg_13_9_inst : DLH_X1 port map( G => N3760, D => N4549, Q => 
                           REGISTERS_13_9_port);
   REGISTERS_reg_13_8_inst : DLH_X1 port map( G => N3760, D => N4547, Q => 
                           REGISTERS_13_8_port);
   REGISTERS_reg_13_7_inst : DLH_X1 port map( G => N3760, D => N4545, Q => 
                           REGISTERS_13_7_port);
   REGISTERS_reg_13_6_inst : DLH_X1 port map( G => N3760, D => N4543, Q => 
                           REGISTERS_13_6_port);
   REGISTERS_reg_13_5_inst : DLH_X1 port map( G => N3760, D => N4541, Q => 
                           REGISTERS_13_5_port);
   REGISTERS_reg_13_4_inst : DLH_X1 port map( G => N3760, D => N4539, Q => 
                           REGISTERS_13_4_port);
   REGISTERS_reg_13_3_inst : DLH_X1 port map( G => N3760, D => N4537, Q => 
                           REGISTERS_13_3_port);
   REGISTERS_reg_13_2_inst : DLH_X1 port map( G => N3760, D => N4535, Q => 
                           REGISTERS_13_2_port);
   REGISTERS_reg_13_1_inst : DLH_X1 port map( G => N3760, D => N4533, Q => 
                           REGISTERS_13_1_port);
   REGISTERS_reg_13_0_inst : DLH_X1 port map( G => N3760, D => N4531, Q => 
                           REGISTERS_13_0_port);
   REGISTERS_reg_14_31_inst : DLH_X1 port map( G => N3696, D => N4593, Q => 
                           REGISTERS_14_31_port);
   REGISTERS_reg_14_30_inst : DLH_X1 port map( G => N3696, D => N4591, Q => 
                           REGISTERS_14_30_port);
   REGISTERS_reg_14_29_inst : DLH_X1 port map( G => N3696, D => N4589, Q => 
                           REGISTERS_14_29_port);
   REGISTERS_reg_14_28_inst : DLH_X1 port map( G => N3696, D => N4587, Q => 
                           REGISTERS_14_28_port);
   REGISTERS_reg_14_27_inst : DLH_X1 port map( G => N3696, D => N4585, Q => 
                           REGISTERS_14_27_port);
   REGISTERS_reg_14_26_inst : DLH_X1 port map( G => N3696, D => N4583, Q => 
                           REGISTERS_14_26_port);
   REGISTERS_reg_14_25_inst : DLH_X1 port map( G => N3696, D => N4581, Q => 
                           REGISTERS_14_25_port);
   REGISTERS_reg_14_24_inst : DLH_X1 port map( G => N3696, D => N4579, Q => 
                           REGISTERS_14_24_port);
   REGISTERS_reg_14_23_inst : DLH_X1 port map( G => N3696, D => N4577, Q => 
                           REGISTERS_14_23_port);
   REGISTERS_reg_14_22_inst : DLH_X1 port map( G => N3696, D => N4575, Q => 
                           REGISTERS_14_22_port);
   REGISTERS_reg_14_21_inst : DLH_X1 port map( G => N3696, D => N4573, Q => 
                           REGISTERS_14_21_port);
   REGISTERS_reg_14_20_inst : DLH_X1 port map( G => N3696, D => N4571, Q => 
                           REGISTERS_14_20_port);
   REGISTERS_reg_14_19_inst : DLH_X1 port map( G => N3696, D => N4569, Q => 
                           REGISTERS_14_19_port);
   REGISTERS_reg_14_18_inst : DLH_X1 port map( G => N3696, D => N4567, Q => 
                           REGISTERS_14_18_port);
   REGISTERS_reg_14_17_inst : DLH_X1 port map( G => N3696, D => N4565, Q => 
                           REGISTERS_14_17_port);
   REGISTERS_reg_14_16_inst : DLH_X1 port map( G => N3696, D => N4563, Q => 
                           REGISTERS_14_16_port);
   REGISTERS_reg_14_15_inst : DLH_X1 port map( G => N3696, D => N4561, Q => 
                           REGISTERS_14_15_port);
   REGISTERS_reg_14_14_inst : DLH_X1 port map( G => N3696, D => N4559, Q => 
                           REGISTERS_14_14_port);
   REGISTERS_reg_14_13_inst : DLH_X1 port map( G => N3696, D => N4557, Q => 
                           REGISTERS_14_13_port);
   REGISTERS_reg_14_12_inst : DLH_X1 port map( G => N3696, D => N4555, Q => 
                           REGISTERS_14_12_port);
   REGISTERS_reg_14_11_inst : DLH_X1 port map( G => N3696, D => N4553, Q => 
                           REGISTERS_14_11_port);
   REGISTERS_reg_14_10_inst : DLH_X1 port map( G => N3696, D => N4551, Q => 
                           REGISTERS_14_10_port);
   REGISTERS_reg_14_9_inst : DLH_X1 port map( G => N3696, D => N4549, Q => 
                           REGISTERS_14_9_port);
   REGISTERS_reg_14_8_inst : DLH_X1 port map( G => N3696, D => N4547, Q => 
                           REGISTERS_14_8_port);
   REGISTERS_reg_14_7_inst : DLH_X1 port map( G => N3696, D => N4545, Q => 
                           REGISTERS_14_7_port);
   REGISTERS_reg_14_6_inst : DLH_X1 port map( G => N3696, D => N4543, Q => 
                           REGISTERS_14_6_port);
   REGISTERS_reg_14_5_inst : DLH_X1 port map( G => N3696, D => N4541, Q => 
                           REGISTERS_14_5_port);
   REGISTERS_reg_14_4_inst : DLH_X1 port map( G => N3696, D => N4539, Q => 
                           REGISTERS_14_4_port);
   REGISTERS_reg_14_3_inst : DLH_X1 port map( G => N3696, D => N4537, Q => 
                           REGISTERS_14_3_port);
   REGISTERS_reg_14_2_inst : DLH_X1 port map( G => N3696, D => N4535, Q => 
                           REGISTERS_14_2_port);
   REGISTERS_reg_14_1_inst : DLH_X1 port map( G => N3696, D => N4533, Q => 
                           REGISTERS_14_1_port);
   REGISTERS_reg_14_0_inst : DLH_X1 port map( G => N3696, D => N4531, Q => 
                           REGISTERS_14_0_port);
   REGISTERS_reg_15_31_inst : DLH_X1 port map( G => N3632, D => N4593, Q => 
                           REGISTERS_15_31_port);
   REGISTERS_reg_15_30_inst : DLH_X1 port map( G => N3632, D => N4591, Q => 
                           REGISTERS_15_30_port);
   REGISTERS_reg_15_29_inst : DLH_X1 port map( G => N3632, D => N4589, Q => 
                           REGISTERS_15_29_port);
   REGISTERS_reg_15_28_inst : DLH_X1 port map( G => N3632, D => N4587, Q => 
                           REGISTERS_15_28_port);
   REGISTERS_reg_15_27_inst : DLH_X1 port map( G => N3632, D => N4585, Q => 
                           REGISTERS_15_27_port);
   REGISTERS_reg_15_26_inst : DLH_X1 port map( G => N3632, D => N4583, Q => 
                           REGISTERS_15_26_port);
   REGISTERS_reg_15_25_inst : DLH_X1 port map( G => N3632, D => N4581, Q => 
                           REGISTERS_15_25_port);
   REGISTERS_reg_15_24_inst : DLH_X1 port map( G => N3632, D => N4579, Q => 
                           REGISTERS_15_24_port);
   REGISTERS_reg_15_23_inst : DLH_X1 port map( G => N3632, D => N4577, Q => 
                           REGISTERS_15_23_port);
   REGISTERS_reg_15_22_inst : DLH_X1 port map( G => N3632, D => N4575, Q => 
                           REGISTERS_15_22_port);
   REGISTERS_reg_15_21_inst : DLH_X1 port map( G => N3632, D => N4573, Q => 
                           REGISTERS_15_21_port);
   REGISTERS_reg_15_20_inst : DLH_X1 port map( G => N3632, D => N4571, Q => 
                           REGISTERS_15_20_port);
   REGISTERS_reg_15_19_inst : DLH_X1 port map( G => N3632, D => N4569, Q => 
                           REGISTERS_15_19_port);
   REGISTERS_reg_15_18_inst : DLH_X1 port map( G => N3632, D => N4567, Q => 
                           REGISTERS_15_18_port);
   REGISTERS_reg_15_17_inst : DLH_X1 port map( G => N3632, D => N4565, Q => 
                           REGISTERS_15_17_port);
   REGISTERS_reg_15_16_inst : DLH_X1 port map( G => N3632, D => N4563, Q => 
                           REGISTERS_15_16_port);
   REGISTERS_reg_15_15_inst : DLH_X1 port map( G => N3632, D => N4561, Q => 
                           REGISTERS_15_15_port);
   REGISTERS_reg_15_14_inst : DLH_X1 port map( G => N3632, D => N4559, Q => 
                           REGISTERS_15_14_port);
   REGISTERS_reg_15_13_inst : DLH_X1 port map( G => N3632, D => N4557, Q => 
                           REGISTERS_15_13_port);
   REGISTERS_reg_15_12_inst : DLH_X1 port map( G => N3632, D => N4555, Q => 
                           REGISTERS_15_12_port);
   REGISTERS_reg_15_11_inst : DLH_X1 port map( G => N3632, D => N4553, Q => 
                           REGISTERS_15_11_port);
   REGISTERS_reg_15_10_inst : DLH_X1 port map( G => N3632, D => N4551, Q => 
                           REGISTERS_15_10_port);
   REGISTERS_reg_15_9_inst : DLH_X1 port map( G => N3632, D => N4549, Q => 
                           REGISTERS_15_9_port);
   REGISTERS_reg_15_8_inst : DLH_X1 port map( G => N3632, D => N4547, Q => 
                           REGISTERS_15_8_port);
   REGISTERS_reg_15_7_inst : DLH_X1 port map( G => N3632, D => N4545, Q => 
                           REGISTERS_15_7_port);
   REGISTERS_reg_15_6_inst : DLH_X1 port map( G => N3632, D => N4543, Q => 
                           REGISTERS_15_6_port);
   REGISTERS_reg_15_5_inst : DLH_X1 port map( G => N3632, D => N4541, Q => 
                           REGISTERS_15_5_port);
   REGISTERS_reg_15_4_inst : DLH_X1 port map( G => N3632, D => N4539, Q => 
                           REGISTERS_15_4_port);
   REGISTERS_reg_15_3_inst : DLH_X1 port map( G => N3632, D => N4537, Q => 
                           REGISTERS_15_3_port);
   REGISTERS_reg_15_2_inst : DLH_X1 port map( G => N3632, D => N4535, Q => 
                           REGISTERS_15_2_port);
   REGISTERS_reg_15_1_inst : DLH_X1 port map( G => N3632, D => N4533, Q => 
                           REGISTERS_15_1_port);
   REGISTERS_reg_15_0_inst : DLH_X1 port map( G => N3632, D => N4531, Q => 
                           REGISTERS_15_0_port);
   REGISTERS_reg_16_31_inst : DLH_X1 port map( G => N3568, D => N4593, Q => 
                           REGISTERS_16_31_port);
   REGISTERS_reg_16_30_inst : DLH_X1 port map( G => N3568, D => N4591, Q => 
                           REGISTERS_16_30_port);
   REGISTERS_reg_16_29_inst : DLH_X1 port map( G => N3568, D => N4589, Q => 
                           REGISTERS_16_29_port);
   REGISTERS_reg_16_28_inst : DLH_X1 port map( G => N3568, D => N4587, Q => 
                           REGISTERS_16_28_port);
   REGISTERS_reg_16_27_inst : DLH_X1 port map( G => N3568, D => N4585, Q => 
                           REGISTERS_16_27_port);
   REGISTERS_reg_16_26_inst : DLH_X1 port map( G => N3568, D => N4583, Q => 
                           REGISTERS_16_26_port);
   REGISTERS_reg_16_25_inst : DLH_X1 port map( G => N3568, D => N4581, Q => 
                           REGISTERS_16_25_port);
   REGISTERS_reg_16_24_inst : DLH_X1 port map( G => N3568, D => N4579, Q => 
                           REGISTERS_16_24_port);
   REGISTERS_reg_16_23_inst : DLH_X1 port map( G => N3568, D => N4577, Q => 
                           REGISTERS_16_23_port);
   REGISTERS_reg_16_22_inst : DLH_X1 port map( G => N3568, D => N4575, Q => 
                           REGISTERS_16_22_port);
   REGISTERS_reg_16_21_inst : DLH_X1 port map( G => N3568, D => N4573, Q => 
                           REGISTERS_16_21_port);
   REGISTERS_reg_16_20_inst : DLH_X1 port map( G => N3568, D => N4571, Q => 
                           REGISTERS_16_20_port);
   REGISTERS_reg_16_19_inst : DLH_X1 port map( G => N3568, D => N4569, Q => 
                           REGISTERS_16_19_port);
   REGISTERS_reg_16_18_inst : DLH_X1 port map( G => N3568, D => N4567, Q => 
                           REGISTERS_16_18_port);
   REGISTERS_reg_16_17_inst : DLH_X1 port map( G => N3568, D => N4565, Q => 
                           REGISTERS_16_17_port);
   REGISTERS_reg_16_16_inst : DLH_X1 port map( G => N3568, D => N4563, Q => 
                           REGISTERS_16_16_port);
   REGISTERS_reg_16_15_inst : DLH_X1 port map( G => N3568, D => N4561, Q => 
                           REGISTERS_16_15_port);
   REGISTERS_reg_16_14_inst : DLH_X1 port map( G => N3568, D => N4559, Q => 
                           REGISTERS_16_14_port);
   REGISTERS_reg_16_13_inst : DLH_X1 port map( G => N3568, D => N4557, Q => 
                           REGISTERS_16_13_port);
   REGISTERS_reg_16_12_inst : DLH_X1 port map( G => N3568, D => N4555, Q => 
                           REGISTERS_16_12_port);
   REGISTERS_reg_16_11_inst : DLH_X1 port map( G => N3568, D => N4553, Q => 
                           REGISTERS_16_11_port);
   REGISTERS_reg_16_10_inst : DLH_X1 port map( G => N3568, D => N4551, Q => 
                           REGISTERS_16_10_port);
   REGISTERS_reg_16_9_inst : DLH_X1 port map( G => N3568, D => N4549, Q => 
                           REGISTERS_16_9_port);
   REGISTERS_reg_16_8_inst : DLH_X1 port map( G => N3568, D => N4547, Q => 
                           REGISTERS_16_8_port);
   REGISTERS_reg_16_7_inst : DLH_X1 port map( G => N3568, D => N4545, Q => 
                           REGISTERS_16_7_port);
   REGISTERS_reg_16_6_inst : DLH_X1 port map( G => N3568, D => N4543, Q => 
                           REGISTERS_16_6_port);
   REGISTERS_reg_16_5_inst : DLH_X1 port map( G => N3568, D => N4541, Q => 
                           REGISTERS_16_5_port);
   REGISTERS_reg_16_4_inst : DLH_X1 port map( G => N3568, D => N4539, Q => 
                           REGISTERS_16_4_port);
   REGISTERS_reg_16_3_inst : DLH_X1 port map( G => N3568, D => N4537, Q => 
                           REGISTERS_16_3_port);
   REGISTERS_reg_16_2_inst : DLH_X1 port map( G => N3568, D => N4535, Q => 
                           REGISTERS_16_2_port);
   REGISTERS_reg_16_1_inst : DLH_X1 port map( G => N3568, D => N4533, Q => 
                           REGISTERS_16_1_port);
   REGISTERS_reg_16_0_inst : DLH_X1 port map( G => N3568, D => N4531, Q => 
                           REGISTERS_16_0_port);
   REGISTERS_reg_17_31_inst : DLH_X1 port map( G => N3504, D => N4593, Q => 
                           REGISTERS_17_31_port);
   REGISTERS_reg_17_30_inst : DLH_X1 port map( G => N3504, D => N4591, Q => 
                           REGISTERS_17_30_port);
   REGISTERS_reg_17_29_inst : DLH_X1 port map( G => N3504, D => N4589, Q => 
                           REGISTERS_17_29_port);
   REGISTERS_reg_17_28_inst : DLH_X1 port map( G => N3504, D => N4587, Q => 
                           REGISTERS_17_28_port);
   REGISTERS_reg_17_27_inst : DLH_X1 port map( G => N3504, D => N4585, Q => 
                           REGISTERS_17_27_port);
   REGISTERS_reg_17_26_inst : DLH_X1 port map( G => N3504, D => N4583, Q => 
                           REGISTERS_17_26_port);
   REGISTERS_reg_17_25_inst : DLH_X1 port map( G => N3504, D => N4581, Q => 
                           REGISTERS_17_25_port);
   REGISTERS_reg_17_24_inst : DLH_X1 port map( G => N3504, D => N4579, Q => 
                           REGISTERS_17_24_port);
   REGISTERS_reg_17_23_inst : DLH_X1 port map( G => N3504, D => N4577, Q => 
                           REGISTERS_17_23_port);
   REGISTERS_reg_17_22_inst : DLH_X1 port map( G => N3504, D => N4575, Q => 
                           REGISTERS_17_22_port);
   REGISTERS_reg_17_21_inst : DLH_X1 port map( G => N3504, D => N4573, Q => 
                           REGISTERS_17_21_port);
   REGISTERS_reg_17_20_inst : DLH_X1 port map( G => N3504, D => N4571, Q => 
                           REGISTERS_17_20_port);
   REGISTERS_reg_17_19_inst : DLH_X1 port map( G => N3504, D => N4569, Q => 
                           REGISTERS_17_19_port);
   REGISTERS_reg_17_18_inst : DLH_X1 port map( G => N3504, D => N4567, Q => 
                           REGISTERS_17_18_port);
   REGISTERS_reg_17_17_inst : DLH_X1 port map( G => N3504, D => N4565, Q => 
                           REGISTERS_17_17_port);
   REGISTERS_reg_17_16_inst : DLH_X1 port map( G => N3504, D => N4563, Q => 
                           REGISTERS_17_16_port);
   REGISTERS_reg_17_15_inst : DLH_X1 port map( G => N3504, D => N4561, Q => 
                           REGISTERS_17_15_port);
   REGISTERS_reg_17_14_inst : DLH_X1 port map( G => N3504, D => N4559, Q => 
                           REGISTERS_17_14_port);
   REGISTERS_reg_17_13_inst : DLH_X1 port map( G => N3504, D => N4557, Q => 
                           REGISTERS_17_13_port);
   REGISTERS_reg_17_12_inst : DLH_X1 port map( G => N3504, D => N4555, Q => 
                           REGISTERS_17_12_port);
   REGISTERS_reg_17_11_inst : DLH_X1 port map( G => N3504, D => N4553, Q => 
                           REGISTERS_17_11_port);
   REGISTERS_reg_17_10_inst : DLH_X1 port map( G => N3504, D => N4551, Q => 
                           REGISTERS_17_10_port);
   REGISTERS_reg_17_9_inst : DLH_X1 port map( G => N3504, D => N4549, Q => 
                           REGISTERS_17_9_port);
   REGISTERS_reg_17_8_inst : DLH_X1 port map( G => N3504, D => N4547, Q => 
                           REGISTERS_17_8_port);
   REGISTERS_reg_17_7_inst : DLH_X1 port map( G => N3504, D => N4545, Q => 
                           REGISTERS_17_7_port);
   REGISTERS_reg_17_6_inst : DLH_X1 port map( G => N3504, D => N4543, Q => 
                           REGISTERS_17_6_port);
   REGISTERS_reg_17_5_inst : DLH_X1 port map( G => N3504, D => N4541, Q => 
                           REGISTERS_17_5_port);
   REGISTERS_reg_17_4_inst : DLH_X1 port map( G => N3504, D => N4539, Q => 
                           REGISTERS_17_4_port);
   REGISTERS_reg_17_3_inst : DLH_X1 port map( G => N3504, D => N4537, Q => 
                           REGISTERS_17_3_port);
   REGISTERS_reg_17_2_inst : DLH_X1 port map( G => N3504, D => N4535, Q => 
                           REGISTERS_17_2_port);
   REGISTERS_reg_17_1_inst : DLH_X1 port map( G => N3504, D => N4533, Q => 
                           REGISTERS_17_1_port);
   REGISTERS_reg_17_0_inst : DLH_X1 port map( G => N3504, D => N4531, Q => 
                           REGISTERS_17_0_port);
   REGISTERS_reg_18_31_inst : DLH_X1 port map( G => N3440, D => N4593, Q => 
                           REGISTERS_18_31_port);
   REGISTERS_reg_18_30_inst : DLH_X1 port map( G => N3440, D => N4591, Q => 
                           REGISTERS_18_30_port);
   REGISTERS_reg_18_29_inst : DLH_X1 port map( G => N3440, D => N4589, Q => 
                           REGISTERS_18_29_port);
   REGISTERS_reg_18_28_inst : DLH_X1 port map( G => N3440, D => N4587, Q => 
                           REGISTERS_18_28_port);
   REGISTERS_reg_18_27_inst : DLH_X1 port map( G => N3440, D => N4585, Q => 
                           REGISTERS_18_27_port);
   REGISTERS_reg_18_26_inst : DLH_X1 port map( G => N3440, D => N4583, Q => 
                           REGISTERS_18_26_port);
   REGISTERS_reg_18_25_inst : DLH_X1 port map( G => N3440, D => N4581, Q => 
                           REGISTERS_18_25_port);
   REGISTERS_reg_18_24_inst : DLH_X1 port map( G => N3440, D => N4579, Q => 
                           REGISTERS_18_24_port);
   REGISTERS_reg_18_23_inst : DLH_X1 port map( G => N3440, D => N4577, Q => 
                           REGISTERS_18_23_port);
   REGISTERS_reg_18_22_inst : DLH_X1 port map( G => N3440, D => N4575, Q => 
                           REGISTERS_18_22_port);
   REGISTERS_reg_18_21_inst : DLH_X1 port map( G => N3440, D => N4573, Q => 
                           REGISTERS_18_21_port);
   REGISTERS_reg_18_20_inst : DLH_X1 port map( G => N3440, D => N4571, Q => 
                           REGISTERS_18_20_port);
   REGISTERS_reg_18_19_inst : DLH_X1 port map( G => N3440, D => N4569, Q => 
                           REGISTERS_18_19_port);
   REGISTERS_reg_18_18_inst : DLH_X1 port map( G => N3440, D => N4567, Q => 
                           REGISTERS_18_18_port);
   REGISTERS_reg_18_17_inst : DLH_X1 port map( G => N3440, D => N4565, Q => 
                           REGISTERS_18_17_port);
   REGISTERS_reg_18_16_inst : DLH_X1 port map( G => N3440, D => N4563, Q => 
                           REGISTERS_18_16_port);
   REGISTERS_reg_18_15_inst : DLH_X1 port map( G => N3440, D => N4561, Q => 
                           REGISTERS_18_15_port);
   REGISTERS_reg_18_14_inst : DLH_X1 port map( G => N3440, D => N4559, Q => 
                           REGISTERS_18_14_port);
   REGISTERS_reg_18_13_inst : DLH_X1 port map( G => N3440, D => N4557, Q => 
                           REGISTERS_18_13_port);
   REGISTERS_reg_18_12_inst : DLH_X1 port map( G => N3440, D => N4555, Q => 
                           REGISTERS_18_12_port);
   REGISTERS_reg_18_11_inst : DLH_X1 port map( G => N3440, D => N4553, Q => 
                           REGISTERS_18_11_port);
   REGISTERS_reg_18_10_inst : DLH_X1 port map( G => N3440, D => N4551, Q => 
                           REGISTERS_18_10_port);
   REGISTERS_reg_18_9_inst : DLH_X1 port map( G => N3440, D => N4549, Q => 
                           REGISTERS_18_9_port);
   REGISTERS_reg_18_8_inst : DLH_X1 port map( G => N3440, D => N4547, Q => 
                           REGISTERS_18_8_port);
   REGISTERS_reg_18_7_inst : DLH_X1 port map( G => N3440, D => N4545, Q => 
                           REGISTERS_18_7_port);
   REGISTERS_reg_18_6_inst : DLH_X1 port map( G => N3440, D => N4543, Q => 
                           REGISTERS_18_6_port);
   REGISTERS_reg_18_5_inst : DLH_X1 port map( G => N3440, D => N4541, Q => 
                           REGISTERS_18_5_port);
   REGISTERS_reg_18_4_inst : DLH_X1 port map( G => N3440, D => N4539, Q => 
                           REGISTERS_18_4_port);
   REGISTERS_reg_18_3_inst : DLH_X1 port map( G => N3440, D => N4537, Q => 
                           REGISTERS_18_3_port);
   REGISTERS_reg_18_2_inst : DLH_X1 port map( G => N3440, D => N4535, Q => 
                           REGISTERS_18_2_port);
   REGISTERS_reg_18_1_inst : DLH_X1 port map( G => N3440, D => N4533, Q => 
                           REGISTERS_18_1_port);
   REGISTERS_reg_18_0_inst : DLH_X1 port map( G => N3440, D => N4531, Q => 
                           REGISTERS_18_0_port);
   REGISTERS_reg_19_31_inst : DLH_X1 port map( G => N3376, D => N4593, Q => 
                           REGISTERS_19_31_port);
   REGISTERS_reg_19_30_inst : DLH_X1 port map( G => N3376, D => N4591, Q => 
                           REGISTERS_19_30_port);
   REGISTERS_reg_19_29_inst : DLH_X1 port map( G => N3376, D => N4589, Q => 
                           REGISTERS_19_29_port);
   REGISTERS_reg_19_28_inst : DLH_X1 port map( G => N3376, D => N4587, Q => 
                           REGISTERS_19_28_port);
   REGISTERS_reg_19_27_inst : DLH_X1 port map( G => N3376, D => N4585, Q => 
                           REGISTERS_19_27_port);
   REGISTERS_reg_19_26_inst : DLH_X1 port map( G => N3376, D => N4583, Q => 
                           REGISTERS_19_26_port);
   REGISTERS_reg_19_25_inst : DLH_X1 port map( G => N3376, D => N4581, Q => 
                           REGISTERS_19_25_port);
   REGISTERS_reg_19_24_inst : DLH_X1 port map( G => N3376, D => N4579, Q => 
                           REGISTERS_19_24_port);
   REGISTERS_reg_19_23_inst : DLH_X1 port map( G => N3376, D => N4577, Q => 
                           REGISTERS_19_23_port);
   REGISTERS_reg_19_22_inst : DLH_X1 port map( G => N3376, D => N4575, Q => 
                           REGISTERS_19_22_port);
   REGISTERS_reg_19_21_inst : DLH_X1 port map( G => N3376, D => N4573, Q => 
                           REGISTERS_19_21_port);
   REGISTERS_reg_19_20_inst : DLH_X1 port map( G => N3376, D => N4571, Q => 
                           REGISTERS_19_20_port);
   REGISTERS_reg_19_19_inst : DLH_X1 port map( G => N3376, D => N4569, Q => 
                           REGISTERS_19_19_port);
   REGISTERS_reg_19_18_inst : DLH_X1 port map( G => N3376, D => N4567, Q => 
                           REGISTERS_19_18_port);
   REGISTERS_reg_19_17_inst : DLH_X1 port map( G => N3376, D => N4565, Q => 
                           REGISTERS_19_17_port);
   REGISTERS_reg_19_16_inst : DLH_X1 port map( G => N3376, D => N4563, Q => 
                           REGISTERS_19_16_port);
   REGISTERS_reg_19_15_inst : DLH_X1 port map( G => N3376, D => N4561, Q => 
                           REGISTERS_19_15_port);
   REGISTERS_reg_19_14_inst : DLH_X1 port map( G => N3376, D => N4559, Q => 
                           REGISTERS_19_14_port);
   REGISTERS_reg_19_13_inst : DLH_X1 port map( G => N3376, D => N4557, Q => 
                           REGISTERS_19_13_port);
   REGISTERS_reg_19_12_inst : DLH_X1 port map( G => N3376, D => N4555, Q => 
                           REGISTERS_19_12_port);
   REGISTERS_reg_19_11_inst : DLH_X1 port map( G => N3376, D => N4553, Q => 
                           REGISTERS_19_11_port);
   REGISTERS_reg_19_10_inst : DLH_X1 port map( G => N3376, D => N4551, Q => 
                           REGISTERS_19_10_port);
   REGISTERS_reg_19_9_inst : DLH_X1 port map( G => N3376, D => N4549, Q => 
                           REGISTERS_19_9_port);
   REGISTERS_reg_19_8_inst : DLH_X1 port map( G => N3376, D => N4547, Q => 
                           REGISTERS_19_8_port);
   REGISTERS_reg_19_7_inst : DLH_X1 port map( G => N3376, D => N4545, Q => 
                           REGISTERS_19_7_port);
   REGISTERS_reg_19_6_inst : DLH_X1 port map( G => N3376, D => N4543, Q => 
                           REGISTERS_19_6_port);
   REGISTERS_reg_19_5_inst : DLH_X1 port map( G => N3376, D => N4541, Q => 
                           REGISTERS_19_5_port);
   REGISTERS_reg_19_4_inst : DLH_X1 port map( G => N3376, D => N4539, Q => 
                           REGISTERS_19_4_port);
   REGISTERS_reg_19_3_inst : DLH_X1 port map( G => N3376, D => N4537, Q => 
                           REGISTERS_19_3_port);
   REGISTERS_reg_19_2_inst : DLH_X1 port map( G => N3376, D => N4535, Q => 
                           REGISTERS_19_2_port);
   REGISTERS_reg_19_1_inst : DLH_X1 port map( G => N3376, D => N4533, Q => 
                           REGISTERS_19_1_port);
   REGISTERS_reg_19_0_inst : DLH_X1 port map( G => N3376, D => N4531, Q => 
                           REGISTERS_19_0_port);
   REGISTERS_reg_20_31_inst : DLH_X1 port map( G => N3312, D => N4593, Q => 
                           REGISTERS_20_31_port);
   REGISTERS_reg_20_30_inst : DLH_X1 port map( G => N3312, D => N4591, Q => 
                           REGISTERS_20_30_port);
   REGISTERS_reg_20_29_inst : DLH_X1 port map( G => N3312, D => N4589, Q => 
                           REGISTERS_20_29_port);
   REGISTERS_reg_20_28_inst : DLH_X1 port map( G => N3312, D => N4587, Q => 
                           REGISTERS_20_28_port);
   REGISTERS_reg_20_27_inst : DLH_X1 port map( G => N3312, D => N4585, Q => 
                           REGISTERS_20_27_port);
   REGISTERS_reg_20_26_inst : DLH_X1 port map( G => N3312, D => N4583, Q => 
                           REGISTERS_20_26_port);
   REGISTERS_reg_20_25_inst : DLH_X1 port map( G => N3312, D => N4581, Q => 
                           REGISTERS_20_25_port);
   REGISTERS_reg_20_24_inst : DLH_X1 port map( G => N3312, D => N4579, Q => 
                           REGISTERS_20_24_port);
   REGISTERS_reg_20_23_inst : DLH_X1 port map( G => N3312, D => N4577, Q => 
                           REGISTERS_20_23_port);
   REGISTERS_reg_20_22_inst : DLH_X1 port map( G => N3312, D => N4575, Q => 
                           REGISTERS_20_22_port);
   REGISTERS_reg_20_21_inst : DLH_X1 port map( G => N3312, D => N4573, Q => 
                           REGISTERS_20_21_port);
   REGISTERS_reg_20_20_inst : DLH_X1 port map( G => N3312, D => N4571, Q => 
                           REGISTERS_20_20_port);
   REGISTERS_reg_20_19_inst : DLH_X1 port map( G => N3312, D => N4569, Q => 
                           REGISTERS_20_19_port);
   REGISTERS_reg_20_18_inst : DLH_X1 port map( G => N3312, D => N4567, Q => 
                           REGISTERS_20_18_port);
   REGISTERS_reg_20_17_inst : DLH_X1 port map( G => N3312, D => N4565, Q => 
                           REGISTERS_20_17_port);
   REGISTERS_reg_20_16_inst : DLH_X1 port map( G => N3312, D => N4563, Q => 
                           REGISTERS_20_16_port);
   REGISTERS_reg_20_15_inst : DLH_X1 port map( G => N3312, D => N4561, Q => 
                           REGISTERS_20_15_port);
   REGISTERS_reg_20_14_inst : DLH_X1 port map( G => N3312, D => N4559, Q => 
                           REGISTERS_20_14_port);
   REGISTERS_reg_20_13_inst : DLH_X1 port map( G => N3312, D => N4557, Q => 
                           REGISTERS_20_13_port);
   REGISTERS_reg_20_12_inst : DLH_X1 port map( G => N3312, D => N4555, Q => 
                           REGISTERS_20_12_port);
   REGISTERS_reg_20_11_inst : DLH_X1 port map( G => N3312, D => N4553, Q => 
                           REGISTERS_20_11_port);
   REGISTERS_reg_20_10_inst : DLH_X1 port map( G => N3312, D => N4551, Q => 
                           REGISTERS_20_10_port);
   REGISTERS_reg_20_9_inst : DLH_X1 port map( G => N3312, D => N4549, Q => 
                           REGISTERS_20_9_port);
   REGISTERS_reg_20_8_inst : DLH_X1 port map( G => N3312, D => N4547, Q => 
                           REGISTERS_20_8_port);
   REGISTERS_reg_20_7_inst : DLH_X1 port map( G => N3312, D => N4545, Q => 
                           REGISTERS_20_7_port);
   REGISTERS_reg_20_6_inst : DLH_X1 port map( G => N3312, D => N4543, Q => 
                           REGISTERS_20_6_port);
   REGISTERS_reg_20_5_inst : DLH_X1 port map( G => N3312, D => N4541, Q => 
                           REGISTERS_20_5_port);
   REGISTERS_reg_20_4_inst : DLH_X1 port map( G => N3312, D => N4539, Q => 
                           REGISTERS_20_4_port);
   REGISTERS_reg_20_3_inst : DLH_X1 port map( G => N3312, D => N4537, Q => 
                           REGISTERS_20_3_port);
   REGISTERS_reg_20_2_inst : DLH_X1 port map( G => N3312, D => N4535, Q => 
                           REGISTERS_20_2_port);
   REGISTERS_reg_20_1_inst : DLH_X1 port map( G => N3312, D => N4533, Q => 
                           REGISTERS_20_1_port);
   REGISTERS_reg_20_0_inst : DLH_X1 port map( G => N3312, D => N4531, Q => 
                           REGISTERS_20_0_port);
   REGISTERS_reg_21_31_inst : DLH_X1 port map( G => N3248, D => N4593, Q => 
                           REGISTERS_21_31_port);
   REGISTERS_reg_21_30_inst : DLH_X1 port map( G => N3248, D => N4591, Q => 
                           REGISTERS_21_30_port);
   REGISTERS_reg_21_29_inst : DLH_X1 port map( G => N3248, D => N4589, Q => 
                           REGISTERS_21_29_port);
   REGISTERS_reg_21_28_inst : DLH_X1 port map( G => N3248, D => N4587, Q => 
                           REGISTERS_21_28_port);
   REGISTERS_reg_21_27_inst : DLH_X1 port map( G => N3248, D => N4585, Q => 
                           REGISTERS_21_27_port);
   REGISTERS_reg_21_26_inst : DLH_X1 port map( G => N3248, D => N4583, Q => 
                           REGISTERS_21_26_port);
   REGISTERS_reg_21_25_inst : DLH_X1 port map( G => N3248, D => N4581, Q => 
                           REGISTERS_21_25_port);
   REGISTERS_reg_21_24_inst : DLH_X1 port map( G => N3248, D => N4579, Q => 
                           REGISTERS_21_24_port);
   REGISTERS_reg_21_23_inst : DLH_X1 port map( G => N3248, D => N4577, Q => 
                           REGISTERS_21_23_port);
   REGISTERS_reg_21_22_inst : DLH_X1 port map( G => N3248, D => N4575, Q => 
                           REGISTERS_21_22_port);
   REGISTERS_reg_21_21_inst : DLH_X1 port map( G => N3248, D => N4573, Q => 
                           REGISTERS_21_21_port);
   REGISTERS_reg_21_20_inst : DLH_X1 port map( G => N3248, D => N4571, Q => 
                           REGISTERS_21_20_port);
   REGISTERS_reg_21_19_inst : DLH_X1 port map( G => N3248, D => N4569, Q => 
                           REGISTERS_21_19_port);
   REGISTERS_reg_21_18_inst : DLH_X1 port map( G => N3248, D => N4567, Q => 
                           REGISTERS_21_18_port);
   REGISTERS_reg_21_17_inst : DLH_X1 port map( G => N3248, D => N4565, Q => 
                           REGISTERS_21_17_port);
   REGISTERS_reg_21_16_inst : DLH_X1 port map( G => N3248, D => N4563, Q => 
                           REGISTERS_21_16_port);
   REGISTERS_reg_21_15_inst : DLH_X1 port map( G => N3248, D => N4561, Q => 
                           REGISTERS_21_15_port);
   REGISTERS_reg_21_14_inst : DLH_X1 port map( G => N3248, D => N4559, Q => 
                           REGISTERS_21_14_port);
   REGISTERS_reg_21_13_inst : DLH_X1 port map( G => N3248, D => N4557, Q => 
                           REGISTERS_21_13_port);
   REGISTERS_reg_21_12_inst : DLH_X1 port map( G => N3248, D => N4555, Q => 
                           REGISTERS_21_12_port);
   REGISTERS_reg_21_11_inst : DLH_X1 port map( G => N3248, D => N4553, Q => 
                           REGISTERS_21_11_port);
   REGISTERS_reg_21_10_inst : DLH_X1 port map( G => N3248, D => N4551, Q => 
                           REGISTERS_21_10_port);
   REGISTERS_reg_21_9_inst : DLH_X1 port map( G => N3248, D => N4549, Q => 
                           REGISTERS_21_9_port);
   REGISTERS_reg_21_8_inst : DLH_X1 port map( G => N3248, D => N4547, Q => 
                           REGISTERS_21_8_port);
   REGISTERS_reg_21_7_inst : DLH_X1 port map( G => N3248, D => N4545, Q => 
                           REGISTERS_21_7_port);
   REGISTERS_reg_21_6_inst : DLH_X1 port map( G => N3248, D => N4543, Q => 
                           REGISTERS_21_6_port);
   REGISTERS_reg_21_5_inst : DLH_X1 port map( G => N3248, D => N4541, Q => 
                           REGISTERS_21_5_port);
   REGISTERS_reg_21_4_inst : DLH_X1 port map( G => N3248, D => N4539, Q => 
                           REGISTERS_21_4_port);
   REGISTERS_reg_21_3_inst : DLH_X1 port map( G => N3248, D => N4537, Q => 
                           REGISTERS_21_3_port);
   REGISTERS_reg_21_2_inst : DLH_X1 port map( G => N3248, D => N4535, Q => 
                           REGISTERS_21_2_port);
   REGISTERS_reg_21_1_inst : DLH_X1 port map( G => N3248, D => N4533, Q => 
                           REGISTERS_21_1_port);
   REGISTERS_reg_21_0_inst : DLH_X1 port map( G => N3248, D => N4531, Q => 
                           REGISTERS_21_0_port);
   REGISTERS_reg_22_31_inst : DLH_X1 port map( G => N3184, D => N4593, Q => 
                           REGISTERS_22_31_port);
   REGISTERS_reg_22_30_inst : DLH_X1 port map( G => N3184, D => N4591, Q => 
                           REGISTERS_22_30_port);
   REGISTERS_reg_22_29_inst : DLH_X1 port map( G => N3184, D => N4589, Q => 
                           REGISTERS_22_29_port);
   REGISTERS_reg_22_28_inst : DLH_X1 port map( G => N3184, D => N4587, Q => 
                           REGISTERS_22_28_port);
   REGISTERS_reg_22_27_inst : DLH_X1 port map( G => N3184, D => N4585, Q => 
                           REGISTERS_22_27_port);
   REGISTERS_reg_22_26_inst : DLH_X1 port map( G => N3184, D => N4583, Q => 
                           REGISTERS_22_26_port);
   REGISTERS_reg_22_25_inst : DLH_X1 port map( G => N3184, D => N4581, Q => 
                           REGISTERS_22_25_port);
   REGISTERS_reg_22_24_inst : DLH_X1 port map( G => N3184, D => N4579, Q => 
                           REGISTERS_22_24_port);
   REGISTERS_reg_22_23_inst : DLH_X1 port map( G => N3184, D => N4577, Q => 
                           REGISTERS_22_23_port);
   REGISTERS_reg_22_22_inst : DLH_X1 port map( G => N3184, D => N4575, Q => 
                           REGISTERS_22_22_port);
   REGISTERS_reg_22_21_inst : DLH_X1 port map( G => N3184, D => N4573, Q => 
                           REGISTERS_22_21_port);
   REGISTERS_reg_22_20_inst : DLH_X1 port map( G => N3184, D => N4571, Q => 
                           REGISTERS_22_20_port);
   REGISTERS_reg_22_19_inst : DLH_X1 port map( G => N3184, D => N4569, Q => 
                           REGISTERS_22_19_port);
   REGISTERS_reg_22_18_inst : DLH_X1 port map( G => N3184, D => N4567, Q => 
                           REGISTERS_22_18_port);
   REGISTERS_reg_22_17_inst : DLH_X1 port map( G => N3184, D => N4565, Q => 
                           REGISTERS_22_17_port);
   REGISTERS_reg_22_16_inst : DLH_X1 port map( G => N3184, D => N4563, Q => 
                           REGISTERS_22_16_port);
   REGISTERS_reg_22_15_inst : DLH_X1 port map( G => N3184, D => N4561, Q => 
                           REGISTERS_22_15_port);
   REGISTERS_reg_22_14_inst : DLH_X1 port map( G => N3184, D => N4559, Q => 
                           REGISTERS_22_14_port);
   REGISTERS_reg_22_13_inst : DLH_X1 port map( G => N3184, D => N4557, Q => 
                           REGISTERS_22_13_port);
   REGISTERS_reg_22_12_inst : DLH_X1 port map( G => N3184, D => N4555, Q => 
                           REGISTERS_22_12_port);
   REGISTERS_reg_22_11_inst : DLH_X1 port map( G => N3184, D => N4553, Q => 
                           REGISTERS_22_11_port);
   REGISTERS_reg_22_10_inst : DLH_X1 port map( G => N3184, D => N4551, Q => 
                           REGISTERS_22_10_port);
   REGISTERS_reg_22_9_inst : DLH_X1 port map( G => N3184, D => N4549, Q => 
                           REGISTERS_22_9_port);
   REGISTERS_reg_22_8_inst : DLH_X1 port map( G => N3184, D => N4547, Q => 
                           REGISTERS_22_8_port);
   REGISTERS_reg_22_7_inst : DLH_X1 port map( G => N3184, D => N4545, Q => 
                           REGISTERS_22_7_port);
   REGISTERS_reg_22_6_inst : DLH_X1 port map( G => N3184, D => N4543, Q => 
                           REGISTERS_22_6_port);
   REGISTERS_reg_22_5_inst : DLH_X1 port map( G => N3184, D => N4541, Q => 
                           REGISTERS_22_5_port);
   REGISTERS_reg_22_4_inst : DLH_X1 port map( G => N3184, D => N4539, Q => 
                           REGISTERS_22_4_port);
   REGISTERS_reg_22_3_inst : DLH_X1 port map( G => N3184, D => N4537, Q => 
                           REGISTERS_22_3_port);
   REGISTERS_reg_22_2_inst : DLH_X1 port map( G => N3184, D => N4535, Q => 
                           REGISTERS_22_2_port);
   REGISTERS_reg_22_1_inst : DLH_X1 port map( G => N3184, D => N4533, Q => 
                           REGISTERS_22_1_port);
   REGISTERS_reg_22_0_inst : DLH_X1 port map( G => N3184, D => N4531, Q => 
                           REGISTERS_22_0_port);
   REGISTERS_reg_23_31_inst : DLH_X1 port map( G => N3120, D => N4593, Q => 
                           REGISTERS_23_31_port);
   REGISTERS_reg_23_30_inst : DLH_X1 port map( G => N3120, D => N4591, Q => 
                           REGISTERS_23_30_port);
   REGISTERS_reg_23_29_inst : DLH_X1 port map( G => N3120, D => N4589, Q => 
                           REGISTERS_23_29_port);
   REGISTERS_reg_23_28_inst : DLH_X1 port map( G => N3120, D => N4587, Q => 
                           REGISTERS_23_28_port);
   REGISTERS_reg_23_27_inst : DLH_X1 port map( G => N3120, D => N4585, Q => 
                           REGISTERS_23_27_port);
   REGISTERS_reg_23_26_inst : DLH_X1 port map( G => N3120, D => N4583, Q => 
                           REGISTERS_23_26_port);
   REGISTERS_reg_23_25_inst : DLH_X1 port map( G => N3120, D => N4581, Q => 
                           REGISTERS_23_25_port);
   REGISTERS_reg_23_24_inst : DLH_X1 port map( G => N3120, D => N4579, Q => 
                           REGISTERS_23_24_port);
   REGISTERS_reg_23_23_inst : DLH_X1 port map( G => N3120, D => N4577, Q => 
                           REGISTERS_23_23_port);
   REGISTERS_reg_23_22_inst : DLH_X1 port map( G => N3120, D => N4575, Q => 
                           REGISTERS_23_22_port);
   REGISTERS_reg_23_21_inst : DLH_X1 port map( G => N3120, D => N4573, Q => 
                           REGISTERS_23_21_port);
   REGISTERS_reg_23_20_inst : DLH_X1 port map( G => N3120, D => N4571, Q => 
                           REGISTERS_23_20_port);
   REGISTERS_reg_23_19_inst : DLH_X1 port map( G => N3120, D => N4569, Q => 
                           REGISTERS_23_19_port);
   REGISTERS_reg_23_18_inst : DLH_X1 port map( G => N3120, D => N4567, Q => 
                           REGISTERS_23_18_port);
   REGISTERS_reg_23_17_inst : DLH_X1 port map( G => N3120, D => N4565, Q => 
                           REGISTERS_23_17_port);
   REGISTERS_reg_23_16_inst : DLH_X1 port map( G => N3120, D => N4563, Q => 
                           REGISTERS_23_16_port);
   REGISTERS_reg_23_15_inst : DLH_X1 port map( G => N3120, D => N4561, Q => 
                           REGISTERS_23_15_port);
   REGISTERS_reg_23_14_inst : DLH_X1 port map( G => N3120, D => N4559, Q => 
                           REGISTERS_23_14_port);
   REGISTERS_reg_23_13_inst : DLH_X1 port map( G => N3120, D => N4557, Q => 
                           REGISTERS_23_13_port);
   REGISTERS_reg_23_12_inst : DLH_X1 port map( G => N3120, D => N4555, Q => 
                           REGISTERS_23_12_port);
   REGISTERS_reg_23_11_inst : DLH_X1 port map( G => N3120, D => N4553, Q => 
                           REGISTERS_23_11_port);
   REGISTERS_reg_23_10_inst : DLH_X1 port map( G => N3120, D => N4551, Q => 
                           REGISTERS_23_10_port);
   REGISTERS_reg_23_9_inst : DLH_X1 port map( G => N3120, D => N4549, Q => 
                           REGISTERS_23_9_port);
   REGISTERS_reg_23_8_inst : DLH_X1 port map( G => N3120, D => N4547, Q => 
                           REGISTERS_23_8_port);
   REGISTERS_reg_23_7_inst : DLH_X1 port map( G => N3120, D => N4545, Q => 
                           REGISTERS_23_7_port);
   REGISTERS_reg_23_6_inst : DLH_X1 port map( G => N3120, D => N4543, Q => 
                           REGISTERS_23_6_port);
   REGISTERS_reg_23_5_inst : DLH_X1 port map( G => N3120, D => N4541, Q => 
                           REGISTERS_23_5_port);
   REGISTERS_reg_23_4_inst : DLH_X1 port map( G => N3120, D => N4539, Q => 
                           REGISTERS_23_4_port);
   REGISTERS_reg_23_3_inst : DLH_X1 port map( G => N3120, D => N4537, Q => 
                           REGISTERS_23_3_port);
   REGISTERS_reg_23_2_inst : DLH_X1 port map( G => N3120, D => N4535, Q => 
                           REGISTERS_23_2_port);
   REGISTERS_reg_23_1_inst : DLH_X1 port map( G => N3120, D => N4533, Q => 
                           REGISTERS_23_1_port);
   REGISTERS_reg_23_0_inst : DLH_X1 port map( G => N3120, D => N4531, Q => 
                           REGISTERS_23_0_port);
   REGISTERS_reg_24_31_inst : DLH_X1 port map( G => N3056, D => N4593, Q => 
                           REGISTERS_24_31_port);
   REGISTERS_reg_24_30_inst : DLH_X1 port map( G => N3056, D => N4591, Q => 
                           REGISTERS_24_30_port);
   REGISTERS_reg_24_29_inst : DLH_X1 port map( G => N3056, D => N4589, Q => 
                           REGISTERS_24_29_port);
   REGISTERS_reg_24_28_inst : DLH_X1 port map( G => N3056, D => N4587, Q => 
                           REGISTERS_24_28_port);
   REGISTERS_reg_24_27_inst : DLH_X1 port map( G => N3056, D => N4585, Q => 
                           REGISTERS_24_27_port);
   REGISTERS_reg_24_26_inst : DLH_X1 port map( G => N3056, D => N4583, Q => 
                           REGISTERS_24_26_port);
   REGISTERS_reg_24_25_inst : DLH_X1 port map( G => N3056, D => N4581, Q => 
                           REGISTERS_24_25_port);
   REGISTERS_reg_24_24_inst : DLH_X1 port map( G => N3056, D => N4579, Q => 
                           REGISTERS_24_24_port);
   REGISTERS_reg_24_23_inst : DLH_X1 port map( G => N3056, D => N4577, Q => 
                           REGISTERS_24_23_port);
   REGISTERS_reg_24_22_inst : DLH_X1 port map( G => N3056, D => N4575, Q => 
                           REGISTERS_24_22_port);
   REGISTERS_reg_24_21_inst : DLH_X1 port map( G => N3056, D => N4573, Q => 
                           REGISTERS_24_21_port);
   REGISTERS_reg_24_20_inst : DLH_X1 port map( G => N3056, D => N4571, Q => 
                           REGISTERS_24_20_port);
   REGISTERS_reg_24_19_inst : DLH_X1 port map( G => N3056, D => N4569, Q => 
                           REGISTERS_24_19_port);
   REGISTERS_reg_24_18_inst : DLH_X1 port map( G => N3056, D => N4567, Q => 
                           REGISTERS_24_18_port);
   REGISTERS_reg_24_17_inst : DLH_X1 port map( G => N3056, D => N4565, Q => 
                           REGISTERS_24_17_port);
   REGISTERS_reg_24_16_inst : DLH_X1 port map( G => N3056, D => N4563, Q => 
                           REGISTERS_24_16_port);
   REGISTERS_reg_24_15_inst : DLH_X1 port map( G => N3056, D => N4561, Q => 
                           REGISTERS_24_15_port);
   REGISTERS_reg_24_14_inst : DLH_X1 port map( G => N3056, D => N4559, Q => 
                           REGISTERS_24_14_port);
   REGISTERS_reg_24_13_inst : DLH_X1 port map( G => N3056, D => N4557, Q => 
                           REGISTERS_24_13_port);
   REGISTERS_reg_24_12_inst : DLH_X1 port map( G => N3056, D => N4555, Q => 
                           REGISTERS_24_12_port);
   REGISTERS_reg_24_11_inst : DLH_X1 port map( G => N3056, D => N4553, Q => 
                           REGISTERS_24_11_port);
   REGISTERS_reg_24_10_inst : DLH_X1 port map( G => N3056, D => N4551, Q => 
                           REGISTERS_24_10_port);
   REGISTERS_reg_24_9_inst : DLH_X1 port map( G => N3056, D => N4549, Q => 
                           REGISTERS_24_9_port);
   REGISTERS_reg_24_8_inst : DLH_X1 port map( G => N3056, D => N4547, Q => 
                           REGISTERS_24_8_port);
   REGISTERS_reg_24_7_inst : DLH_X1 port map( G => N3056, D => N4545, Q => 
                           REGISTERS_24_7_port);
   REGISTERS_reg_24_6_inst : DLH_X1 port map( G => N3056, D => N4543, Q => 
                           REGISTERS_24_6_port);
   REGISTERS_reg_24_5_inst : DLH_X1 port map( G => N3056, D => N4541, Q => 
                           REGISTERS_24_5_port);
   REGISTERS_reg_24_4_inst : DLH_X1 port map( G => N3056, D => N4539, Q => 
                           REGISTERS_24_4_port);
   REGISTERS_reg_24_3_inst : DLH_X1 port map( G => N3056, D => N4537, Q => 
                           REGISTERS_24_3_port);
   REGISTERS_reg_24_2_inst : DLH_X1 port map( G => N3056, D => N4535, Q => 
                           REGISTERS_24_2_port);
   REGISTERS_reg_24_1_inst : DLH_X1 port map( G => N3056, D => N4533, Q => 
                           REGISTERS_24_1_port);
   REGISTERS_reg_24_0_inst : DLH_X1 port map( G => N3056, D => N4531, Q => 
                           REGISTERS_24_0_port);
   REGISTERS_reg_25_31_inst : DLH_X1 port map( G => N2992, D => N4593, Q => 
                           REGISTERS_25_31_port);
   REGISTERS_reg_25_30_inst : DLH_X1 port map( G => N2992, D => N4591, Q => 
                           REGISTERS_25_30_port);
   REGISTERS_reg_25_29_inst : DLH_X1 port map( G => N2992, D => N4589, Q => 
                           REGISTERS_25_29_port);
   REGISTERS_reg_25_28_inst : DLH_X1 port map( G => N2992, D => N4587, Q => 
                           REGISTERS_25_28_port);
   REGISTERS_reg_25_27_inst : DLH_X1 port map( G => N2992, D => N4585, Q => 
                           REGISTERS_25_27_port);
   REGISTERS_reg_25_26_inst : DLH_X1 port map( G => N2992, D => N4583, Q => 
                           REGISTERS_25_26_port);
   REGISTERS_reg_25_25_inst : DLH_X1 port map( G => N2992, D => N4581, Q => 
                           REGISTERS_25_25_port);
   REGISTERS_reg_25_24_inst : DLH_X1 port map( G => N2992, D => N4579, Q => 
                           REGISTERS_25_24_port);
   REGISTERS_reg_25_23_inst : DLH_X1 port map( G => N2992, D => N4577, Q => 
                           REGISTERS_25_23_port);
   REGISTERS_reg_25_22_inst : DLH_X1 port map( G => N2992, D => N4575, Q => 
                           REGISTERS_25_22_port);
   REGISTERS_reg_25_21_inst : DLH_X1 port map( G => N2992, D => N4573, Q => 
                           REGISTERS_25_21_port);
   REGISTERS_reg_25_20_inst : DLH_X1 port map( G => N2992, D => N4571, Q => 
                           REGISTERS_25_20_port);
   REGISTERS_reg_25_19_inst : DLH_X1 port map( G => N2992, D => N4569, Q => 
                           REGISTERS_25_19_port);
   REGISTERS_reg_25_18_inst : DLH_X1 port map( G => N2992, D => N4567, Q => 
                           REGISTERS_25_18_port);
   REGISTERS_reg_25_17_inst : DLH_X1 port map( G => N2992, D => N4565, Q => 
                           REGISTERS_25_17_port);
   REGISTERS_reg_25_16_inst : DLH_X1 port map( G => N2992, D => N4563, Q => 
                           REGISTERS_25_16_port);
   REGISTERS_reg_25_15_inst : DLH_X1 port map( G => N2992, D => N4561, Q => 
                           REGISTERS_25_15_port);
   REGISTERS_reg_25_14_inst : DLH_X1 port map( G => N2992, D => N4559, Q => 
                           REGISTERS_25_14_port);
   REGISTERS_reg_25_13_inst : DLH_X1 port map( G => N2992, D => N4557, Q => 
                           REGISTERS_25_13_port);
   REGISTERS_reg_25_12_inst : DLH_X1 port map( G => N2992, D => N4555, Q => 
                           REGISTERS_25_12_port);
   REGISTERS_reg_25_11_inst : DLH_X1 port map( G => N2992, D => N4553, Q => 
                           REGISTERS_25_11_port);
   REGISTERS_reg_25_10_inst : DLH_X1 port map( G => N2992, D => N4551, Q => 
                           REGISTERS_25_10_port);
   REGISTERS_reg_25_9_inst : DLH_X1 port map( G => N2992, D => N4549, Q => 
                           REGISTERS_25_9_port);
   REGISTERS_reg_25_8_inst : DLH_X1 port map( G => N2992, D => N4547, Q => 
                           REGISTERS_25_8_port);
   REGISTERS_reg_25_7_inst : DLH_X1 port map( G => N2992, D => N4545, Q => 
                           REGISTERS_25_7_port);
   REGISTERS_reg_25_6_inst : DLH_X1 port map( G => N2992, D => N4543, Q => 
                           REGISTERS_25_6_port);
   REGISTERS_reg_25_5_inst : DLH_X1 port map( G => N2992, D => N4541, Q => 
                           REGISTERS_25_5_port);
   REGISTERS_reg_25_4_inst : DLH_X1 port map( G => N2992, D => N4539, Q => 
                           REGISTERS_25_4_port);
   REGISTERS_reg_25_3_inst : DLH_X1 port map( G => N2992, D => N4537, Q => 
                           REGISTERS_25_3_port);
   REGISTERS_reg_25_2_inst : DLH_X1 port map( G => N2992, D => N4535, Q => 
                           REGISTERS_25_2_port);
   REGISTERS_reg_25_1_inst : DLH_X1 port map( G => N2992, D => N4533, Q => 
                           REGISTERS_25_1_port);
   REGISTERS_reg_25_0_inst : DLH_X1 port map( G => N2992, D => N4531, Q => 
                           REGISTERS_25_0_port);
   REGISTERS_reg_26_31_inst : DLH_X1 port map( G => N2928, D => N4593, Q => 
                           REGISTERS_26_31_port);
   REGISTERS_reg_26_30_inst : DLH_X1 port map( G => N2928, D => N4591, Q => 
                           REGISTERS_26_30_port);
   REGISTERS_reg_26_29_inst : DLH_X1 port map( G => N2928, D => N4589, Q => 
                           REGISTERS_26_29_port);
   REGISTERS_reg_26_28_inst : DLH_X1 port map( G => N2928, D => N4587, Q => 
                           REGISTERS_26_28_port);
   REGISTERS_reg_26_27_inst : DLH_X1 port map( G => N2928, D => N4585, Q => 
                           REGISTERS_26_27_port);
   REGISTERS_reg_26_26_inst : DLH_X1 port map( G => N2928, D => N4583, Q => 
                           REGISTERS_26_26_port);
   REGISTERS_reg_26_25_inst : DLH_X1 port map( G => N2928, D => N4581, Q => 
                           REGISTERS_26_25_port);
   REGISTERS_reg_26_24_inst : DLH_X1 port map( G => N2928, D => N4579, Q => 
                           REGISTERS_26_24_port);
   REGISTERS_reg_26_23_inst : DLH_X1 port map( G => N2928, D => N4577, Q => 
                           REGISTERS_26_23_port);
   REGISTERS_reg_26_22_inst : DLH_X1 port map( G => N2928, D => N4575, Q => 
                           REGISTERS_26_22_port);
   REGISTERS_reg_26_21_inst : DLH_X1 port map( G => N2928, D => N4573, Q => 
                           REGISTERS_26_21_port);
   REGISTERS_reg_26_20_inst : DLH_X1 port map( G => N2928, D => N4571, Q => 
                           REGISTERS_26_20_port);
   REGISTERS_reg_26_19_inst : DLH_X1 port map( G => N2928, D => N4569, Q => 
                           REGISTERS_26_19_port);
   REGISTERS_reg_26_18_inst : DLH_X1 port map( G => N2928, D => N4567, Q => 
                           REGISTERS_26_18_port);
   REGISTERS_reg_26_17_inst : DLH_X1 port map( G => N2928, D => N4565, Q => 
                           REGISTERS_26_17_port);
   REGISTERS_reg_26_16_inst : DLH_X1 port map( G => N2928, D => N4563, Q => 
                           REGISTERS_26_16_port);
   REGISTERS_reg_26_15_inst : DLH_X1 port map( G => N2928, D => N4561, Q => 
                           REGISTERS_26_15_port);
   REGISTERS_reg_26_14_inst : DLH_X1 port map( G => N2928, D => N4559, Q => 
                           REGISTERS_26_14_port);
   REGISTERS_reg_26_13_inst : DLH_X1 port map( G => N2928, D => N4557, Q => 
                           REGISTERS_26_13_port);
   REGISTERS_reg_26_12_inst : DLH_X1 port map( G => N2928, D => N4555, Q => 
                           REGISTERS_26_12_port);
   REGISTERS_reg_26_11_inst : DLH_X1 port map( G => N2928, D => N4553, Q => 
                           REGISTERS_26_11_port);
   REGISTERS_reg_26_10_inst : DLH_X1 port map( G => N2928, D => N4551, Q => 
                           REGISTERS_26_10_port);
   REGISTERS_reg_26_9_inst : DLH_X1 port map( G => N2928, D => N4549, Q => 
                           REGISTERS_26_9_port);
   REGISTERS_reg_26_8_inst : DLH_X1 port map( G => N2928, D => N4547, Q => 
                           REGISTERS_26_8_port);
   REGISTERS_reg_26_7_inst : DLH_X1 port map( G => N2928, D => N4545, Q => 
                           REGISTERS_26_7_port);
   REGISTERS_reg_26_6_inst : DLH_X1 port map( G => N2928, D => N4543, Q => 
                           REGISTERS_26_6_port);
   REGISTERS_reg_26_5_inst : DLH_X1 port map( G => N2928, D => N4541, Q => 
                           REGISTERS_26_5_port);
   REGISTERS_reg_26_4_inst : DLH_X1 port map( G => N2928, D => N4539, Q => 
                           REGISTERS_26_4_port);
   REGISTERS_reg_26_3_inst : DLH_X1 port map( G => N2928, D => N4537, Q => 
                           REGISTERS_26_3_port);
   REGISTERS_reg_26_2_inst : DLH_X1 port map( G => N2928, D => N4535, Q => 
                           REGISTERS_26_2_port);
   REGISTERS_reg_26_1_inst : DLH_X1 port map( G => N2928, D => N4533, Q => 
                           REGISTERS_26_1_port);
   REGISTERS_reg_26_0_inst : DLH_X1 port map( G => N2928, D => N4531, Q => 
                           REGISTERS_26_0_port);
   REGISTERS_reg_27_31_inst : DLH_X1 port map( G => N2864, D => N4593, Q => 
                           REGISTERS_27_31_port);
   REGISTERS_reg_27_30_inst : DLH_X1 port map( G => N2864, D => N4591, Q => 
                           REGISTERS_27_30_port);
   REGISTERS_reg_27_29_inst : DLH_X1 port map( G => N2864, D => N4589, Q => 
                           REGISTERS_27_29_port);
   REGISTERS_reg_27_28_inst : DLH_X1 port map( G => N2864, D => N4587, Q => 
                           REGISTERS_27_28_port);
   REGISTERS_reg_27_27_inst : DLH_X1 port map( G => N2864, D => N4585, Q => 
                           REGISTERS_27_27_port);
   REGISTERS_reg_27_26_inst : DLH_X1 port map( G => N2864, D => N4583, Q => 
                           REGISTERS_27_26_port);
   REGISTERS_reg_27_25_inst : DLH_X1 port map( G => N2864, D => N4581, Q => 
                           REGISTERS_27_25_port);
   REGISTERS_reg_27_24_inst : DLH_X1 port map( G => N2864, D => N4579, Q => 
                           REGISTERS_27_24_port);
   REGISTERS_reg_27_23_inst : DLH_X1 port map( G => N2864, D => N4577, Q => 
                           REGISTERS_27_23_port);
   REGISTERS_reg_27_22_inst : DLH_X1 port map( G => N2864, D => N4575, Q => 
                           REGISTERS_27_22_port);
   REGISTERS_reg_27_21_inst : DLH_X1 port map( G => N2864, D => N4573, Q => 
                           REGISTERS_27_21_port);
   REGISTERS_reg_27_20_inst : DLH_X1 port map( G => N2864, D => N4571, Q => 
                           REGISTERS_27_20_port);
   REGISTERS_reg_27_19_inst : DLH_X1 port map( G => N2864, D => N4569, Q => 
                           REGISTERS_27_19_port);
   REGISTERS_reg_27_18_inst : DLH_X1 port map( G => N2864, D => N4567, Q => 
                           REGISTERS_27_18_port);
   REGISTERS_reg_27_17_inst : DLH_X1 port map( G => N2864, D => N4565, Q => 
                           REGISTERS_27_17_port);
   REGISTERS_reg_27_16_inst : DLH_X1 port map( G => N2864, D => N4563, Q => 
                           REGISTERS_27_16_port);
   REGISTERS_reg_27_15_inst : DLH_X1 port map( G => N2864, D => N4561, Q => 
                           REGISTERS_27_15_port);
   REGISTERS_reg_27_14_inst : DLH_X1 port map( G => N2864, D => N4559, Q => 
                           REGISTERS_27_14_port);
   REGISTERS_reg_27_13_inst : DLH_X1 port map( G => N2864, D => N4557, Q => 
                           REGISTERS_27_13_port);
   REGISTERS_reg_27_12_inst : DLH_X1 port map( G => N2864, D => N4555, Q => 
                           REGISTERS_27_12_port);
   REGISTERS_reg_27_11_inst : DLH_X1 port map( G => N2864, D => N4553, Q => 
                           REGISTERS_27_11_port);
   REGISTERS_reg_27_10_inst : DLH_X1 port map( G => N2864, D => N4551, Q => 
                           REGISTERS_27_10_port);
   REGISTERS_reg_27_9_inst : DLH_X1 port map( G => N2864, D => N4549, Q => 
                           REGISTERS_27_9_port);
   REGISTERS_reg_27_8_inst : DLH_X1 port map( G => N2864, D => N4547, Q => 
                           REGISTERS_27_8_port);
   REGISTERS_reg_27_7_inst : DLH_X1 port map( G => N2864, D => N4545, Q => 
                           REGISTERS_27_7_port);
   REGISTERS_reg_27_6_inst : DLH_X1 port map( G => N2864, D => N4543, Q => 
                           REGISTERS_27_6_port);
   REGISTERS_reg_27_5_inst : DLH_X1 port map( G => N2864, D => N4541, Q => 
                           REGISTERS_27_5_port);
   REGISTERS_reg_27_4_inst : DLH_X1 port map( G => N2864, D => N4539, Q => 
                           REGISTERS_27_4_port);
   REGISTERS_reg_27_3_inst : DLH_X1 port map( G => N2864, D => N4537, Q => 
                           REGISTERS_27_3_port);
   REGISTERS_reg_27_2_inst : DLH_X1 port map( G => N2864, D => N4535, Q => 
                           REGISTERS_27_2_port);
   REGISTERS_reg_27_1_inst : DLH_X1 port map( G => N2864, D => N4533, Q => 
                           REGISTERS_27_1_port);
   REGISTERS_reg_27_0_inst : DLH_X1 port map( G => N2864, D => N4531, Q => 
                           REGISTERS_27_0_port);
   REGISTERS_reg_28_31_inst : DLH_X1 port map( G => N2800, D => N4593, Q => 
                           REGISTERS_28_31_port);
   REGISTERS_reg_28_30_inst : DLH_X1 port map( G => N2800, D => N4591, Q => 
                           REGISTERS_28_30_port);
   REGISTERS_reg_28_29_inst : DLH_X1 port map( G => N2800, D => N4589, Q => 
                           REGISTERS_28_29_port);
   REGISTERS_reg_28_28_inst : DLH_X1 port map( G => N2800, D => N4587, Q => 
                           REGISTERS_28_28_port);
   REGISTERS_reg_28_27_inst : DLH_X1 port map( G => N2800, D => N4585, Q => 
                           REGISTERS_28_27_port);
   REGISTERS_reg_28_26_inst : DLH_X1 port map( G => N2800, D => N4583, Q => 
                           REGISTERS_28_26_port);
   REGISTERS_reg_28_25_inst : DLH_X1 port map( G => N2800, D => N4581, Q => 
                           REGISTERS_28_25_port);
   REGISTERS_reg_28_24_inst : DLH_X1 port map( G => N2800, D => N4579, Q => 
                           REGISTERS_28_24_port);
   REGISTERS_reg_28_23_inst : DLH_X1 port map( G => N2800, D => N4577, Q => 
                           REGISTERS_28_23_port);
   REGISTERS_reg_28_22_inst : DLH_X1 port map( G => N2800, D => N4575, Q => 
                           REGISTERS_28_22_port);
   REGISTERS_reg_28_21_inst : DLH_X1 port map( G => N2800, D => N4573, Q => 
                           REGISTERS_28_21_port);
   REGISTERS_reg_28_20_inst : DLH_X1 port map( G => N2800, D => N4571, Q => 
                           REGISTERS_28_20_port);
   REGISTERS_reg_28_19_inst : DLH_X1 port map( G => N2800, D => N4569, Q => 
                           REGISTERS_28_19_port);
   REGISTERS_reg_28_18_inst : DLH_X1 port map( G => N2800, D => N4567, Q => 
                           REGISTERS_28_18_port);
   REGISTERS_reg_28_17_inst : DLH_X1 port map( G => N2800, D => N4565, Q => 
                           REGISTERS_28_17_port);
   REGISTERS_reg_28_16_inst : DLH_X1 port map( G => N2800, D => N4563, Q => 
                           REGISTERS_28_16_port);
   REGISTERS_reg_28_15_inst : DLH_X1 port map( G => N2800, D => N4561, Q => 
                           REGISTERS_28_15_port);
   REGISTERS_reg_28_14_inst : DLH_X1 port map( G => N2800, D => N4559, Q => 
                           REGISTERS_28_14_port);
   REGISTERS_reg_28_13_inst : DLH_X1 port map( G => N2800, D => N4557, Q => 
                           REGISTERS_28_13_port);
   REGISTERS_reg_28_12_inst : DLH_X1 port map( G => N2800, D => N4555, Q => 
                           REGISTERS_28_12_port);
   REGISTERS_reg_28_11_inst : DLH_X1 port map( G => N2800, D => N4553, Q => 
                           REGISTERS_28_11_port);
   REGISTERS_reg_28_10_inst : DLH_X1 port map( G => N2800, D => N4551, Q => 
                           REGISTERS_28_10_port);
   REGISTERS_reg_28_9_inst : DLH_X1 port map( G => N2800, D => N4549, Q => 
                           REGISTERS_28_9_port);
   REGISTERS_reg_28_8_inst : DLH_X1 port map( G => N2800, D => N4547, Q => 
                           REGISTERS_28_8_port);
   REGISTERS_reg_28_7_inst : DLH_X1 port map( G => N2800, D => N4545, Q => 
                           REGISTERS_28_7_port);
   REGISTERS_reg_28_6_inst : DLH_X1 port map( G => N2800, D => N4543, Q => 
                           REGISTERS_28_6_port);
   REGISTERS_reg_28_5_inst : DLH_X1 port map( G => N2800, D => N4541, Q => 
                           REGISTERS_28_5_port);
   REGISTERS_reg_28_4_inst : DLH_X1 port map( G => N2800, D => N4539, Q => 
                           REGISTERS_28_4_port);
   REGISTERS_reg_28_3_inst : DLH_X1 port map( G => N2800, D => N4537, Q => 
                           REGISTERS_28_3_port);
   REGISTERS_reg_28_2_inst : DLH_X1 port map( G => N2800, D => N4535, Q => 
                           REGISTERS_28_2_port);
   REGISTERS_reg_28_1_inst : DLH_X1 port map( G => N2800, D => N4533, Q => 
                           REGISTERS_28_1_port);
   REGISTERS_reg_28_0_inst : DLH_X1 port map( G => N2800, D => N4531, Q => 
                           REGISTERS_28_0_port);
   REGISTERS_reg_29_31_inst : DLH_X1 port map( G => N2736, D => N4593, Q => 
                           REGISTERS_29_31_port);
   REGISTERS_reg_29_30_inst : DLH_X1 port map( G => N2736, D => N4591, Q => 
                           REGISTERS_29_30_port);
   REGISTERS_reg_29_29_inst : DLH_X1 port map( G => N2736, D => N4589, Q => 
                           REGISTERS_29_29_port);
   REGISTERS_reg_29_28_inst : DLH_X1 port map( G => N2736, D => N4587, Q => 
                           REGISTERS_29_28_port);
   REGISTERS_reg_29_27_inst : DLH_X1 port map( G => N2736, D => N4585, Q => 
                           REGISTERS_29_27_port);
   REGISTERS_reg_29_26_inst : DLH_X1 port map( G => N2736, D => N4583, Q => 
                           REGISTERS_29_26_port);
   REGISTERS_reg_29_25_inst : DLH_X1 port map( G => N2736, D => N4581, Q => 
                           REGISTERS_29_25_port);
   REGISTERS_reg_29_24_inst : DLH_X1 port map( G => N2736, D => N4579, Q => 
                           REGISTERS_29_24_port);
   REGISTERS_reg_29_23_inst : DLH_X1 port map( G => N2736, D => N4577, Q => 
                           REGISTERS_29_23_port);
   REGISTERS_reg_29_22_inst : DLH_X1 port map( G => N2736, D => N4575, Q => 
                           REGISTERS_29_22_port);
   REGISTERS_reg_29_21_inst : DLH_X1 port map( G => N2736, D => N4573, Q => 
                           REGISTERS_29_21_port);
   REGISTERS_reg_29_20_inst : DLH_X1 port map( G => N2736, D => N4571, Q => 
                           REGISTERS_29_20_port);
   REGISTERS_reg_29_19_inst : DLH_X1 port map( G => N2736, D => N4569, Q => 
                           REGISTERS_29_19_port);
   REGISTERS_reg_29_18_inst : DLH_X1 port map( G => N2736, D => N4567, Q => 
                           REGISTERS_29_18_port);
   REGISTERS_reg_29_17_inst : DLH_X1 port map( G => N2736, D => N4565, Q => 
                           REGISTERS_29_17_port);
   REGISTERS_reg_29_16_inst : DLH_X1 port map( G => N2736, D => N4563, Q => 
                           REGISTERS_29_16_port);
   REGISTERS_reg_29_15_inst : DLH_X1 port map( G => N2736, D => N4561, Q => 
                           REGISTERS_29_15_port);
   REGISTERS_reg_29_14_inst : DLH_X1 port map( G => N2736, D => N4559, Q => 
                           REGISTERS_29_14_port);
   REGISTERS_reg_29_13_inst : DLH_X1 port map( G => N2736, D => N4557, Q => 
                           REGISTERS_29_13_port);
   REGISTERS_reg_29_12_inst : DLH_X1 port map( G => N2736, D => N4555, Q => 
                           REGISTERS_29_12_port);
   REGISTERS_reg_29_11_inst : DLH_X1 port map( G => N2736, D => N4553, Q => 
                           REGISTERS_29_11_port);
   REGISTERS_reg_29_10_inst : DLH_X1 port map( G => N2736, D => N4551, Q => 
                           REGISTERS_29_10_port);
   REGISTERS_reg_29_9_inst : DLH_X1 port map( G => N2736, D => N4549, Q => 
                           REGISTERS_29_9_port);
   REGISTERS_reg_29_8_inst : DLH_X1 port map( G => N2736, D => N4547, Q => 
                           REGISTERS_29_8_port);
   REGISTERS_reg_29_7_inst : DLH_X1 port map( G => N2736, D => N4545, Q => 
                           REGISTERS_29_7_port);
   REGISTERS_reg_29_6_inst : DLH_X1 port map( G => N2736, D => N4543, Q => 
                           REGISTERS_29_6_port);
   REGISTERS_reg_29_5_inst : DLH_X1 port map( G => N2736, D => N4541, Q => 
                           REGISTERS_29_5_port);
   REGISTERS_reg_29_4_inst : DLH_X1 port map( G => N2736, D => N4539, Q => 
                           REGISTERS_29_4_port);
   REGISTERS_reg_29_3_inst : DLH_X1 port map( G => N2736, D => N4537, Q => 
                           REGISTERS_29_3_port);
   REGISTERS_reg_29_2_inst : DLH_X1 port map( G => N2736, D => N4535, Q => 
                           REGISTERS_29_2_port);
   REGISTERS_reg_29_1_inst : DLH_X1 port map( G => N2736, D => N4533, Q => 
                           REGISTERS_29_1_port);
   REGISTERS_reg_29_0_inst : DLH_X1 port map( G => N2736, D => N4531, Q => 
                           REGISTERS_29_0_port);
   REGISTERS_reg_30_31_inst : DLH_X1 port map( G => N2672, D => N4593, Q => 
                           REGISTERS_30_31_port);
   REGISTERS_reg_30_30_inst : DLH_X1 port map( G => N2672, D => N4591, Q => 
                           REGISTERS_30_30_port);
   REGISTERS_reg_30_29_inst : DLH_X1 port map( G => N2672, D => N4589, Q => 
                           REGISTERS_30_29_port);
   REGISTERS_reg_30_28_inst : DLH_X1 port map( G => N2672, D => N4587, Q => 
                           REGISTERS_30_28_port);
   REGISTERS_reg_30_27_inst : DLH_X1 port map( G => N2672, D => N4585, Q => 
                           REGISTERS_30_27_port);
   REGISTERS_reg_30_26_inst : DLH_X1 port map( G => N2672, D => N4583, Q => 
                           REGISTERS_30_26_port);
   REGISTERS_reg_30_25_inst : DLH_X1 port map( G => N2672, D => N4581, Q => 
                           REGISTERS_30_25_port);
   REGISTERS_reg_30_24_inst : DLH_X1 port map( G => N2672, D => N4579, Q => 
                           REGISTERS_30_24_port);
   REGISTERS_reg_30_23_inst : DLH_X1 port map( G => N2672, D => N4577, Q => 
                           REGISTERS_30_23_port);
   REGISTERS_reg_30_22_inst : DLH_X1 port map( G => N2672, D => N4575, Q => 
                           REGISTERS_30_22_port);
   REGISTERS_reg_30_21_inst : DLH_X1 port map( G => N2672, D => N4573, Q => 
                           REGISTERS_30_21_port);
   REGISTERS_reg_30_20_inst : DLH_X1 port map( G => N2672, D => N4571, Q => 
                           REGISTERS_30_20_port);
   REGISTERS_reg_30_19_inst : DLH_X1 port map( G => N2672, D => N4569, Q => 
                           REGISTERS_30_19_port);
   REGISTERS_reg_30_18_inst : DLH_X1 port map( G => N2672, D => N4567, Q => 
                           REGISTERS_30_18_port);
   REGISTERS_reg_30_17_inst : DLH_X1 port map( G => N2672, D => N4565, Q => 
                           REGISTERS_30_17_port);
   REGISTERS_reg_30_16_inst : DLH_X1 port map( G => N2672, D => N4563, Q => 
                           REGISTERS_30_16_port);
   REGISTERS_reg_30_15_inst : DLH_X1 port map( G => N2672, D => N4561, Q => 
                           REGISTERS_30_15_port);
   REGISTERS_reg_30_14_inst : DLH_X1 port map( G => N2672, D => N4559, Q => 
                           REGISTERS_30_14_port);
   REGISTERS_reg_30_13_inst : DLH_X1 port map( G => N2672, D => N4557, Q => 
                           REGISTERS_30_13_port);
   REGISTERS_reg_30_12_inst : DLH_X1 port map( G => N2672, D => N4555, Q => 
                           REGISTERS_30_12_port);
   REGISTERS_reg_30_11_inst : DLH_X1 port map( G => N2672, D => N4553, Q => 
                           REGISTERS_30_11_port);
   REGISTERS_reg_30_10_inst : DLH_X1 port map( G => N2672, D => N4551, Q => 
                           REGISTERS_30_10_port);
   REGISTERS_reg_30_9_inst : DLH_X1 port map( G => N2672, D => N4549, Q => 
                           REGISTERS_30_9_port);
   REGISTERS_reg_30_8_inst : DLH_X1 port map( G => N2672, D => N4547, Q => 
                           REGISTERS_30_8_port);
   REGISTERS_reg_30_7_inst : DLH_X1 port map( G => N2672, D => N4545, Q => 
                           REGISTERS_30_7_port);
   REGISTERS_reg_30_6_inst : DLH_X1 port map( G => N2672, D => N4543, Q => 
                           REGISTERS_30_6_port);
   REGISTERS_reg_30_5_inst : DLH_X1 port map( G => N2672, D => N4541, Q => 
                           REGISTERS_30_5_port);
   REGISTERS_reg_30_4_inst : DLH_X1 port map( G => N2672, D => N4539, Q => 
                           REGISTERS_30_4_port);
   REGISTERS_reg_30_3_inst : DLH_X1 port map( G => N2672, D => N4537, Q => 
                           REGISTERS_30_3_port);
   REGISTERS_reg_30_2_inst : DLH_X1 port map( G => N2672, D => N4535, Q => 
                           REGISTERS_30_2_port);
   REGISTERS_reg_30_1_inst : DLH_X1 port map( G => N2672, D => N4533, Q => 
                           REGISTERS_30_1_port);
   REGISTERS_reg_30_0_inst : DLH_X1 port map( G => N2672, D => N4531, Q => 
                           REGISTERS_30_0_port);
   REGISTERS_reg_31_31_inst : DLH_X1 port map( G => N2608, D => N4593, Q => 
                           REGISTERS_31_31_port);
   REGISTERS_reg_31_30_inst : DLH_X1 port map( G => N2608, D => N4591, Q => 
                           REGISTERS_31_30_port);
   REGISTERS_reg_31_29_inst : DLH_X1 port map( G => N2608, D => N4589, Q => 
                           REGISTERS_31_29_port);
   REGISTERS_reg_31_28_inst : DLH_X1 port map( G => N2608, D => N4587, Q => 
                           REGISTERS_31_28_port);
   REGISTERS_reg_31_27_inst : DLH_X1 port map( G => N2608, D => N4585, Q => 
                           REGISTERS_31_27_port);
   REGISTERS_reg_31_26_inst : DLH_X1 port map( G => N2608, D => N4583, Q => 
                           REGISTERS_31_26_port);
   REGISTERS_reg_31_25_inst : DLH_X1 port map( G => N2608, D => N4581, Q => 
                           REGISTERS_31_25_port);
   REGISTERS_reg_31_24_inst : DLH_X1 port map( G => N2608, D => N4579, Q => 
                           REGISTERS_31_24_port);
   REGISTERS_reg_31_23_inst : DLH_X1 port map( G => N2608, D => N4577, Q => 
                           REGISTERS_31_23_port);
   REGISTERS_reg_31_22_inst : DLH_X1 port map( G => N2608, D => N4575, Q => 
                           REGISTERS_31_22_port);
   REGISTERS_reg_31_21_inst : DLH_X1 port map( G => N2608, D => N4573, Q => 
                           REGISTERS_31_21_port);
   REGISTERS_reg_31_20_inst : DLH_X1 port map( G => N2608, D => N4571, Q => 
                           REGISTERS_31_20_port);
   REGISTERS_reg_31_19_inst : DLH_X1 port map( G => N2608, D => N4569, Q => 
                           REGISTERS_31_19_port);
   REGISTERS_reg_31_18_inst : DLH_X1 port map( G => N2608, D => N4567, Q => 
                           REGISTERS_31_18_port);
   REGISTERS_reg_31_17_inst : DLH_X1 port map( G => N2608, D => N4565, Q => 
                           REGISTERS_31_17_port);
   REGISTERS_reg_31_16_inst : DLH_X1 port map( G => N2608, D => N4563, Q => 
                           REGISTERS_31_16_port);
   REGISTERS_reg_31_15_inst : DLH_X1 port map( G => N2608, D => N4561, Q => 
                           REGISTERS_31_15_port);
   REGISTERS_reg_31_14_inst : DLH_X1 port map( G => N2608, D => N4559, Q => 
                           REGISTERS_31_14_port);
   REGISTERS_reg_31_13_inst : DLH_X1 port map( G => N2608, D => N4557, Q => 
                           REGISTERS_31_13_port);
   REGISTERS_reg_31_12_inst : DLH_X1 port map( G => N2608, D => N4555, Q => 
                           REGISTERS_31_12_port);
   REGISTERS_reg_31_11_inst : DLH_X1 port map( G => N2608, D => N4553, Q => 
                           REGISTERS_31_11_port);
   REGISTERS_reg_31_10_inst : DLH_X1 port map( G => N2608, D => N4551, Q => 
                           REGISTERS_31_10_port);
   REGISTERS_reg_31_9_inst : DLH_X1 port map( G => N2608, D => N4549, Q => 
                           REGISTERS_31_9_port);
   REGISTERS_reg_31_8_inst : DLH_X1 port map( G => N2608, D => N4547, Q => 
                           REGISTERS_31_8_port);
   REGISTERS_reg_31_7_inst : DLH_X1 port map( G => N2608, D => N4545, Q => 
                           REGISTERS_31_7_port);
   REGISTERS_reg_31_6_inst : DLH_X1 port map( G => N2608, D => N4543, Q => 
                           REGISTERS_31_6_port);
   REGISTERS_reg_31_5_inst : DLH_X1 port map( G => N2608, D => N4541, Q => 
                           REGISTERS_31_5_port);
   REGISTERS_reg_31_4_inst : DLH_X1 port map( G => N2608, D => N4539, Q => 
                           REGISTERS_31_4_port);
   REGISTERS_reg_31_3_inst : DLH_X1 port map( G => N2608, D => N4537, Q => 
                           REGISTERS_31_3_port);
   REGISTERS_reg_31_2_inst : DLH_X1 port map( G => N2608, D => N4535, Q => 
                           REGISTERS_31_2_port);
   REGISTERS_reg_31_1_inst : DLH_X1 port map( G => N2608, D => N4533, Q => 
                           REGISTERS_31_1_port);
   REGISTERS_reg_31_0_inst : DLH_X1 port map( G => N2608, D => N4531, Q => 
                           REGISTERS_31_0_port);
   OUT1_reg_31_inst : DLH_X1 port map( G => N2480, D => N2481, Q => OUT1(31));
   OUT1_reg_30_inst : DLH_X1 port map( G => N2480, D => N2479, Q => OUT1(30));
   OUT1_reg_29_inst : DLH_X1 port map( G => N2480, D => N2477, Q => OUT1(29));
   OUT1_reg_28_inst : DLH_X1 port map( G => N2480, D => N2475, Q => OUT1(28));
   OUT1_reg_27_inst : DLH_X1 port map( G => N2480, D => N2473, Q => OUT1(27));
   OUT1_reg_26_inst : DLH_X1 port map( G => N2480, D => N2471, Q => OUT1(26));
   OUT1_reg_25_inst : DLH_X1 port map( G => N2480, D => N2469, Q => OUT1(25));
   OUT1_reg_24_inst : DLH_X1 port map( G => N2480, D => N2467, Q => OUT1(24));
   OUT1_reg_23_inst : DLH_X1 port map( G => N2480, D => N2465, Q => OUT1(23));
   OUT1_reg_22_inst : DLH_X1 port map( G => N2480, D => N2463, Q => OUT1(22));
   OUT1_reg_21_inst : DLH_X1 port map( G => N2480, D => N2461, Q => OUT1(21));
   OUT1_reg_20_inst : DLH_X1 port map( G => N2480, D => N2459, Q => OUT1(20));
   OUT1_reg_19_inst : DLH_X1 port map( G => N2480, D => N2457, Q => OUT1(19));
   OUT1_reg_18_inst : DLH_X1 port map( G => N2480, D => N2455, Q => OUT1(18));
   OUT1_reg_17_inst : DLH_X1 port map( G => N2480, D => N2453, Q => OUT1(17));
   OUT1_reg_16_inst : DLH_X1 port map( G => N2480, D => N2451, Q => OUT1(16));
   OUT1_reg_15_inst : DLH_X1 port map( G => N2480, D => N2449, Q => OUT1(15));
   OUT1_reg_14_inst : DLH_X1 port map( G => N2480, D => N2447, Q => OUT1(14));
   OUT1_reg_13_inst : DLH_X1 port map( G => N2480, D => N2445, Q => OUT1(13));
   OUT1_reg_12_inst : DLH_X1 port map( G => N2480, D => N2443, Q => OUT1(12));
   OUT1_reg_11_inst : DLH_X1 port map( G => N2480, D => N2441, Q => OUT1(11));
   OUT1_reg_10_inst : DLH_X1 port map( G => N2480, D => N2439, Q => OUT1(10));
   OUT1_reg_9_inst : DLH_X1 port map( G => N2480, D => N2437, Q => OUT1(9));
   OUT1_reg_8_inst : DLH_X1 port map( G => N2480, D => N2435, Q => OUT1(8));
   OUT1_reg_7_inst : DLH_X1 port map( G => N2480, D => N2433, Q => OUT1(7));
   OUT1_reg_6_inst : DLH_X1 port map( G => N2480, D => N2431, Q => OUT1(6));
   OUT1_reg_5_inst : DLH_X1 port map( G => N2480, D => N2429, Q => OUT1(5));
   OUT1_reg_4_inst : DLH_X1 port map( G => N2480, D => N2427, Q => OUT1(4));
   OUT1_reg_3_inst : DLH_X1 port map( G => N2480, D => N2425, Q => OUT1(3));
   OUT1_reg_2_inst : DLH_X1 port map( G => N2480, D => N2423, Q => OUT1(2));
   OUT1_reg_1_inst : DLH_X1 port map( G => N2480, D => N2421, Q => OUT1(1));
   OUT1_reg_0_inst : DLH_X1 port map( G => N2480, D => N2419, Q => OUT1(0));
   OUT2_reg_31_inst : DLH_X1 port map( G => N2544, D => N2545, Q => OUT2(31));
   OUT2_reg_30_inst : DLH_X1 port map( G => N2544, D => N2543, Q => OUT2(30));
   OUT2_reg_29_inst : DLH_X1 port map( G => N2544, D => N2541, Q => OUT2(29));
   OUT2_reg_28_inst : DLH_X1 port map( G => N2544, D => N2539, Q => OUT2(28));
   OUT2_reg_27_inst : DLH_X1 port map( G => N2544, D => N2537, Q => OUT2(27));
   OUT2_reg_26_inst : DLH_X1 port map( G => N2544, D => N2535, Q => OUT2(26));
   OUT2_reg_25_inst : DLH_X1 port map( G => N2544, D => N2533, Q => OUT2(25));
   OUT2_reg_24_inst : DLH_X1 port map( G => N2544, D => N2531, Q => OUT2(24));
   OUT2_reg_23_inst : DLH_X1 port map( G => N2544, D => N2529, Q => OUT2(23));
   OUT2_reg_22_inst : DLH_X1 port map( G => N2544, D => N2527, Q => OUT2(22));
   OUT2_reg_21_inst : DLH_X1 port map( G => N2544, D => N2525, Q => OUT2(21));
   OUT2_reg_20_inst : DLH_X1 port map( G => N2544, D => N2523, Q => OUT2(20));
   OUT2_reg_19_inst : DLH_X1 port map( G => N2544, D => N2521, Q => OUT2(19));
   OUT2_reg_18_inst : DLH_X1 port map( G => N2544, D => N2519, Q => OUT2(18));
   OUT2_reg_17_inst : DLH_X1 port map( G => N2544, D => N2517, Q => OUT2(17));
   OUT2_reg_16_inst : DLH_X1 port map( G => N2544, D => N2515, Q => OUT2(16));
   OUT2_reg_15_inst : DLH_X1 port map( G => N2544, D => N2513, Q => OUT2(15));
   OUT2_reg_14_inst : DLH_X1 port map( G => N2544, D => N2511, Q => OUT2(14));
   OUT2_reg_13_inst : DLH_X1 port map( G => N2544, D => N2509, Q => OUT2(13));
   OUT2_reg_12_inst : DLH_X1 port map( G => N2544, D => N2507, Q => OUT2(12));
   OUT2_reg_11_inst : DLH_X1 port map( G => N2544, D => N2505, Q => OUT2(11));
   OUT2_reg_10_inst : DLH_X1 port map( G => N2544, D => N2503, Q => OUT2(10));
   OUT2_reg_9_inst : DLH_X1 port map( G => N2544, D => N2501, Q => OUT2(9));
   OUT2_reg_8_inst : DLH_X1 port map( G => N2544, D => N2499, Q => OUT2(8));
   OUT2_reg_7_inst : DLH_X1 port map( G => N2544, D => N2497, Q => OUT2(7));
   OUT2_reg_6_inst : DLH_X1 port map( G => N2544, D => N2495, Q => OUT2(6));
   OUT2_reg_5_inst : DLH_X1 port map( G => N2544, D => N2493, Q => OUT2(5));
   OUT2_reg_4_inst : DLH_X1 port map( G => N2544, D => N2491, Q => OUT2(4));
   OUT2_reg_3_inst : DLH_X1 port map( G => N2544, D => N2489, Q => OUT2(3));
   OUT2_reg_2_inst : DLH_X1 port map( G => N2544, D => N2487, Q => OUT2(2));
   OUT2_reg_1_inst : DLH_X1 port map( G => N2544, D => N2485, Q => OUT2(1));
   OUT2_reg_0_inst : DLH_X1 port map( G => N2544, D => N2483, Q => OUT2(0));
   U3 : OAI21_X4 port map( B1 => n2, B2 => n14, A => RESET, ZN => N3568);
   U4 : OAI21_X4 port map( B1 => n9, B2 => n13, A => RESET, ZN => N3632);
   U5 : OAI21_X4 port map( B1 => n3, B2 => n14, A => RESET, ZN => N3504);
   U6 : OAI21_X4 port map( B1 => n8, B2 => n13, A => RESET, ZN => N3696);
   U7 : OAI21_X4 port map( B1 => n4, B2 => n14, A => RESET, ZN => N3440);
   U8 : OAI21_X4 port map( B1 => n7, B2 => n13, A => RESET, ZN => N3760);
   U9 : OAI21_X4 port map( B1 => n5, B2 => n14, A => RESET, ZN => N3376);
   U10 : OAI21_X4 port map( B1 => n6, B2 => n13, A => RESET, ZN => N3824);
   U11 : OAI21_X4 port map( B1 => n6, B2 => n14, A => RESET, ZN => N3312);
   U12 : OAI21_X4 port map( B1 => n5, B2 => n13, A => RESET, ZN => N3888);
   U13 : OAI21_X4 port map( B1 => n7, B2 => n14, A => RESET, ZN => N3248);
   U14 : OAI21_X4 port map( B1 => n4, B2 => n13, A => RESET, ZN => N3952);
   U15 : OAI21_X4 port map( B1 => n8, B2 => n14, A => RESET, ZN => N3184);
   U16 : OAI21_X4 port map( B1 => n3, B2 => n13, A => RESET, ZN => N4016);
   U17 : OAI21_X4 port map( B1 => n9, B2 => n14, A => RESET, ZN => N3120);
   U18 : OAI21_X4 port map( B1 => n2, B2 => n13, A => RESET, ZN => N4080);
   U19 : OAI21_X4 port map( B1 => n1, B2 => n9, A => RESET, ZN => N4144);
   U20 : OAI21_X4 port map( B1 => n2, B2 => n15, A => RESET, ZN => N3056);
   U21 : OAI21_X4 port map( B1 => n3, B2 => n15, A => RESET, ZN => N2992);
   U22 : OAI21_X4 port map( B1 => n1, B2 => n8, A => RESET, ZN => N4208);
   U23 : OAI21_X4 port map( B1 => n1, B2 => n7, A => RESET, ZN => N4272);
   U24 : OAI21_X4 port map( B1 => n4, B2 => n15, A => RESET, ZN => N2928);
   U25 : OAI21_X4 port map( B1 => n5, B2 => n15, A => RESET, ZN => N2864);
   U26 : OAI21_X4 port map( B1 => n1, B2 => n6, A => RESET, ZN => N4336);
   U27 : OAI21_X4 port map( B1 => n1, B2 => n5, A => RESET, ZN => N4400);
   U28 : OAI21_X4 port map( B1 => n6, B2 => n15, A => RESET, ZN => N2800);
   U29 : OAI21_X4 port map( B1 => n7, B2 => n15, A => RESET, ZN => N2736);
   U30 : OAI21_X4 port map( B1 => n1, B2 => n4, A => RESET, ZN => N4464);
   U31 : OAI21_X4 port map( B1 => n1, B2 => n3, A => RESET, ZN => N4528);
   U32 : OAI21_X4 port map( B1 => n8, B2 => n15, A => RESET, ZN => N2672);
   U33 : OAI21_X4 port map( B1 => n9, B2 => n15, A => RESET, ZN => N2608);
   U34 : OAI21_X4 port map( B1 => n1, B2 => n2, A => RESET, ZN => N4592);
   U35 : AND2_X2 port map( A1 => n1771, A2 => n1754, ZN => n1190);
   U36 : NAND2_X2 port map( A1 => n1141, A2 => n1118, ZN => n59);
   U37 : AND2_X2 port map( A1 => n1753, A2 => n1754, ZN => n1166);
   U38 : NAND2_X2 port map( A1 => n1115, A2 => n1118, ZN => n27);
   U39 : NAND2_X2 port map( A1 => n1775, A2 => n1756, ZN => n1197);
   U40 : AND2_X2 port map( A1 => n1149, A2 => n1116, ZN => n77);
   U41 : AND2_X2 port map( A1 => n1775, A2 => n1758, ZN => n1205);
   U42 : AND2_X2 port map( A1 => n1754, A2 => n1762, ZN => n1176);
   U43 : NAND2_X2 port map( A1 => n1149, A2 => n1123, ZN => n80);
   U44 : NAND2_X2 port map( A1 => n1118, A2 => n1128, ZN => n41);
   U45 : NAND2_X2 port map( A1 => n1771, A2 => n1759, ZN => n1192);
   U46 : NAND2_X2 port map( A1 => n1753, A2 => n1756, ZN => n1163);
   U47 : AND2_X2 port map( A1 => n1141, A2 => n1122, ZN => n70);
   U48 : AND2_X2 port map( A1 => n1115, A2 => n1116, ZN => n31);
   U49 : AND2_X2 port map( A1 => n1771, A2 => n1758, ZN => n1195);
   U50 : AND2_X2 port map( A1 => n1753, A2 => n1758, ZN => n1171);
   U51 : NOR3_X2 port map( A1 => ADD_RD1(1), A2 => ADD_RD1(2), A3 => n85, ZN =>
                           n1758);
   U52 : NAND2_X2 port map( A1 => n1128, A2 => n1123, ZN => n48);
   U53 : NAND2_X2 port map( A1 => n1775, A2 => n1759, ZN => n1202);
   U54 : NAND2_X2 port map( A1 => n1756, A2 => n1762, ZN => n1173);
   U55 : AND2_X2 port map( A1 => n1141, A2 => n1116, ZN => n63);
   U56 : AND2_X2 port map( A1 => n1149, A2 => n1122, ZN => n84);
   U57 : AND2_X2 port map( A1 => n1115, A2 => n1122, ZN => n38);
   U58 : NOR3_X2 port map( A1 => ADD_RD2(1), A2 => ADD_RD2(2), A3 => n85, ZN =>
                           n1122);
   U59 : AND2_X2 port map( A1 => n1775, A2 => n1754, ZN => n1200);
   U60 : AND2_X2 port map( A1 => n1758, A2 => n1762, ZN => n1181);
   U61 : NAND2_X2 port map( A1 => n1149, A2 => n1118, ZN => n73);
   U62 : NAND2_X2 port map( A1 => n1115, A2 => n1123, ZN => n34);
   U63 : NAND2_X2 port map( A1 => n1753, A2 => n1759, ZN => n1168);
   U64 : NAND2_X2 port map( A1 => n1771, A2 => n1756, ZN => n1187);
   U65 : AND2_X2 port map( A1 => n1122, A2 => n1128, ZN => n52);
   U66 : AND2_X2 port map( A1 => n1142, A2 => n1116, ZN => n62);
   U67 : NAND2_X2 port map( A1 => n1141, A2 => n1123, ZN => n66);
   U68 : NAND2_X2 port map( A1 => n1755, A2 => n1759, ZN => n1167);
   U69 : NAND2_X2 port map( A1 => n1756, A2 => n1763, ZN => n1172);
   U70 : AND2_X2 port map( A1 => n1772, A2 => n1758, ZN => n1194);
   U71 : AND2_X2 port map( A1 => n1776, A2 => n1754, ZN => n1199);
   U72 : AND2_X2 port map( A1 => n1117, A2 => n1122, ZN => n37);
   U73 : AND2_X2 port map( A1 => n1116, A2 => n1129, ZN => n44);
   U74 : NAND2_X2 port map( A1 => n1150, A2 => n1118, ZN => n71);
   U75 : NAND2_X2 port map( A1 => n1755, A2 => n1756, ZN => n1162);
   U76 : NAND2_X2 port map( A1 => n1763, A2 => n1759, ZN => n1177);
   U77 : AND2_X2 port map( A1 => n1772, A2 => n1754, ZN => n1189);
   U78 : AND2_X2 port map( A1 => n1776, A2 => n1758, ZN => n1204);
   U79 : AND2_X2 port map( A1 => n1117, A2 => n1116, ZN => n30);
   U80 : AND2_X2 port map( A1 => n1122, A2 => n1129, ZN => n51);
   U81 : NAND2_X2 port map( A1 => n1142, A2 => n1118, ZN => n57);
   U82 : NAND2_X2 port map( A1 => n1150, A2 => n1123, ZN => n78);
   U83 : NAND2_X2 port map( A1 => n1772, A2 => n1759, ZN => n1191);
   U84 : NAND2_X2 port map( A1 => n1776, A2 => n1756, ZN => n1196);
   U85 : AND2_X2 port map( A1 => n1755, A2 => n1758, ZN => n1170);
   U86 : AND2_X2 port map( A1 => n1754, A2 => n1763, ZN => n1175);
   U87 : AND2_X2 port map( A1 => n1142, A2 => n1122, ZN => n69);
   U88 : AND2_X2 port map( A1 => n1150, A2 => n1116, ZN => n76);
   U89 : NAND2_X2 port map( A1 => n1117, A2 => n1123, ZN => n32);
   U90 : NAND2_X2 port map( A1 => n1118, A2 => n1129, ZN => n39);
   U91 : NAND2_X2 port map( A1 => n1762, A2 => n1759, ZN => n1178);
   U92 : AND2_X2 port map( A1 => n1116, A2 => n1128, ZN => n45);
   U93 : NAND2_X2 port map( A1 => n1776, A2 => n1759, ZN => n1201);
   U94 : NOR3_X2 port map( A1 => n85, A2 => ADD_RD1(2), A3 => n1777, ZN => 
                           n1759);
   U95 : NAND2_X2 port map( A1 => n1772, A2 => n1756, ZN => n1186);
   U96 : AND2_X2 port map( A1 => n1755, A2 => n1754, ZN => n1165);
   U97 : AND2_X2 port map( A1 => n1758, A2 => n1763, ZN => n1180);
   U98 : AND2_X2 port map( A1 => n1150, A2 => n1122, ZN => n83);
   U99 : NAND2_X2 port map( A1 => n1117, A2 => n1118, ZN => n25);
   U100 : NAND2_X2 port map( A1 => n1129, A2 => n1123, ZN => n46);
   U101 : NAND2_X2 port map( A1 => n1142, A2 => n1123, ZN => n64);
   U102 : NOR3_X2 port map( A1 => n85, A2 => ADD_RD2(2), A3 => n1152, ZN => 
                           n1123);
   U103 : AND2_X1 port map( A1 => RESET, A2 => DATAIN(31), ZN => N4593);
   U104 : AND2_X1 port map( A1 => DATAIN(30), A2 => RESET, ZN => N4591);
   U105 : AND2_X1 port map( A1 => DATAIN(29), A2 => RESET, ZN => N4589);
   U106 : AND2_X1 port map( A1 => DATAIN(28), A2 => RESET, ZN => N4587);
   U107 : AND2_X1 port map( A1 => DATAIN(27), A2 => RESET, ZN => N4585);
   U108 : AND2_X1 port map( A1 => DATAIN(26), A2 => RESET, ZN => N4583);
   U109 : AND2_X1 port map( A1 => DATAIN(25), A2 => RESET, ZN => N4581);
   U110 : AND2_X1 port map( A1 => DATAIN(24), A2 => RESET, ZN => N4579);
   U111 : AND2_X1 port map( A1 => DATAIN(23), A2 => RESET, ZN => N4577);
   U112 : AND2_X1 port map( A1 => DATAIN(22), A2 => RESET, ZN => N4575);
   U113 : AND2_X1 port map( A1 => DATAIN(21), A2 => RESET, ZN => N4573);
   U114 : AND2_X1 port map( A1 => DATAIN(20), A2 => RESET, ZN => N4571);
   U115 : AND2_X1 port map( A1 => DATAIN(19), A2 => RESET, ZN => N4569);
   U116 : AND2_X1 port map( A1 => DATAIN(18), A2 => RESET, ZN => N4567);
   U117 : AND2_X1 port map( A1 => DATAIN(17), A2 => RESET, ZN => N4565);
   U118 : AND2_X1 port map( A1 => DATAIN(16), A2 => RESET, ZN => N4563);
   U119 : AND2_X1 port map( A1 => DATAIN(15), A2 => RESET, ZN => N4561);
   U120 : AND2_X1 port map( A1 => DATAIN(14), A2 => RESET, ZN => N4559);
   U121 : AND2_X1 port map( A1 => DATAIN(13), A2 => RESET, ZN => N4557);
   U122 : AND2_X1 port map( A1 => DATAIN(12), A2 => RESET, ZN => N4555);
   U123 : AND2_X1 port map( A1 => DATAIN(11), A2 => RESET, ZN => N4553);
   U124 : AND2_X1 port map( A1 => DATAIN(10), A2 => RESET, ZN => N4551);
   U125 : AND2_X1 port map( A1 => DATAIN(9), A2 => RESET, ZN => N4549);
   U126 : AND2_X1 port map( A1 => DATAIN(8), A2 => RESET, ZN => N4547);
   U127 : AND2_X1 port map( A1 => DATAIN(7), A2 => RESET, ZN => N4545);
   U128 : AND2_X1 port map( A1 => DATAIN(6), A2 => RESET, ZN => N4543);
   U129 : AND2_X1 port map( A1 => DATAIN(5), A2 => RESET, ZN => N4541);
   U130 : AND2_X1 port map( A1 => DATAIN(4), A2 => RESET, ZN => N4539);
   U131 : AND2_X1 port map( A1 => DATAIN(3), A2 => RESET, ZN => N4537);
   U132 : AND2_X1 port map( A1 => DATAIN(2), A2 => RESET, ZN => N4535);
   U133 : AND2_X1 port map( A1 => DATAIN(1), A2 => RESET, ZN => N4533);
   U134 : AND2_X1 port map( A1 => DATAIN(0), A2 => RESET, ZN => N4531);
   U135 : NAND3_X1 port map( A1 => n10, A2 => n11, A3 => n12, ZN => n1);
   U136 : NAND3_X1 port map( A1 => n12, A2 => n11, A3 => ADD_WR(3), ZN => n13);
   U137 : INV_X1 port map( A => ADD_WR(4), ZN => n11);
   U138 : NAND3_X1 port map( A1 => n12, A2 => n10, A3 => ADD_WR(4), ZN => n14);
   U139 : INV_X1 port map( A => ADD_WR(3), ZN => n10);
   U140 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => n18, ZN => n2);
   U141 : NAND3_X1 port map( A1 => n16, A2 => n17, A3 => ADD_WR(0), ZN => n3);
   U142 : NAND3_X1 port map( A1 => n18, A2 => n17, A3 => ADD_WR(1), ZN => n4);
   U143 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n17, A3 => ADD_WR(1), ZN =>
                           n5);
   U144 : INV_X1 port map( A => ADD_WR(2), ZN => n17);
   U145 : NAND3_X1 port map( A1 => n18, A2 => n16, A3 => ADD_WR(2), ZN => n6);
   U146 : NAND3_X1 port map( A1 => ADD_WR(0), A2 => n16, A3 => ADD_WR(2), ZN =>
                           n7);
   U147 : INV_X1 port map( A => ADD_WR(1), ZN => n16);
   U148 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => n18, A3 => ADD_WR(2), ZN =>
                           n8);
   U149 : INV_X1 port map( A => ADD_WR(0), ZN => n18);
   U150 : NAND3_X1 port map( A1 => ADD_WR(3), A2 => n12, A3 => ADD_WR(4), ZN =>
                           n15);
   U151 : AND2_X1 port map( A1 => WR, A2 => ENABLE, ZN => n12);
   U152 : NAND3_X1 port map( A1 => ADD_WR(1), A2 => ADD_WR(0), A3 => ADD_WR(2),
                           ZN => n9);
   U153 : NAND2_X1 port map( A1 => n19, A2 => n20, ZN => N2545);
   U154 : NOR4_X1 port map( A1 => n21, A2 => n22, A3 => n23, A4 => n24, ZN => 
                           n20);
   U155 : OAI221_X1 port map( B1 => n25, B2 => n26, C1 => n27, C2 => n28, A => 
                           n29, ZN => n24);
   U156 : AOI22_X1 port map( A1 => REGISTERS_28_31_port, A2 => n30, B1 => 
                           REGISTERS_29_31_port, B2 => n31, ZN => n29);
   U157 : OAI221_X1 port map( B1 => n32, B2 => n33, C1 => n34, C2 => n35, A => 
                           n36, ZN => n23);
   U158 : AOI22_X1 port map( A1 => REGISTERS_24_31_port, A2 => n37, B1 => 
                           REGISTERS_25_31_port, B2 => n38, ZN => n36);
   U159 : OAI221_X1 port map( B1 => n39, B2 => n40, C1 => n41, C2 => n42, A => 
                           n43, ZN => n22);
   U160 : AOI22_X1 port map( A1 => REGISTERS_20_31_port, A2 => n44, B1 => 
                           REGISTERS_21_31_port, B2 => n45, ZN => n43);
   U161 : OAI221_X1 port map( B1 => n46, B2 => n47, C1 => n48, C2 => n49, A => 
                           n50, ZN => n21);
   U162 : AOI22_X1 port map( A1 => REGISTERS_16_31_port, A2 => n51, B1 => 
                           REGISTERS_17_31_port, B2 => n52, ZN => n50);
   U163 : NOR4_X1 port map( A1 => n53, A2 => n54, A3 => n55, A4 => n56, ZN => 
                           n19);
   U164 : OAI221_X1 port map( B1 => n57, B2 => n58, C1 => n59, C2 => n60, A => 
                           n61, ZN => n56);
   U165 : AOI22_X1 port map( A1 => REGISTERS_12_31_port, A2 => n62, B1 => 
                           REGISTERS_13_31_port, B2 => n63, ZN => n61);
   U166 : OAI221_X1 port map( B1 => n64, B2 => n65, C1 => n66, C2 => n67, A => 
                           n68, ZN => n55);
   U167 : AOI22_X1 port map( A1 => REGISTERS_8_31_port, A2 => n69, B1 => 
                           REGISTERS_9_31_port, B2 => n70, ZN => n68);
   U168 : OAI221_X1 port map( B1 => n71, B2 => n72, C1 => n73, C2 => n74, A => 
                           n75, ZN => n54);
   U169 : AOI22_X1 port map( A1 => REGISTERS_4_31_port, A2 => n76, B1 => 
                           REGISTERS_5_31_port, B2 => n77, ZN => n75);
   U170 : OAI221_X1 port map( B1 => n78, B2 => n79, C1 => n80, C2 => n81, A => 
                           n82, ZN => n53);
   U171 : AOI22_X1 port map( A1 => REGISTERS_0_31_port, A2 => n83, B1 => 
                           REGISTERS_1_31_port, B2 => n84, ZN => n82);
   U172 : OR2_X1 port map( A1 => RD2, A2 => n85, ZN => N2544);
   U173 : NAND2_X1 port map( A1 => n86, A2 => n87, ZN => N2543);
   U174 : NOR4_X1 port map( A1 => n88, A2 => n89, A3 => n90, A4 => n91, ZN => 
                           n87);
   U175 : OAI221_X1 port map( B1 => n25, B2 => n92, C1 => n27, C2 => n93, A => 
                           n94, ZN => n91);
   U176 : AOI22_X1 port map( A1 => REGISTERS_28_30_port, A2 => n30, B1 => 
                           REGISTERS_29_30_port, B2 => n31, ZN => n94);
   U177 : OAI221_X1 port map( B1 => n32, B2 => n95, C1 => n34, C2 => n96, A => 
                           n97, ZN => n90);
   U178 : AOI22_X1 port map( A1 => REGISTERS_24_30_port, A2 => n37, B1 => 
                           REGISTERS_25_30_port, B2 => n38, ZN => n97);
   U179 : OAI221_X1 port map( B1 => n39, B2 => n98, C1 => n41, C2 => n99, A => 
                           n100, ZN => n89);
   U180 : AOI22_X1 port map( A1 => REGISTERS_20_30_port, A2 => n44, B1 => 
                           REGISTERS_21_30_port, B2 => n45, ZN => n100);
   U181 : OAI221_X1 port map( B1 => n46, B2 => n101, C1 => n48, C2 => n102, A 
                           => n103, ZN => n88);
   U182 : AOI22_X1 port map( A1 => REGISTERS_16_30_port, A2 => n51, B1 => 
                           REGISTERS_17_30_port, B2 => n52, ZN => n103);
   U183 : NOR4_X1 port map( A1 => n104, A2 => n105, A3 => n106, A4 => n107, ZN 
                           => n86);
   U184 : OAI221_X1 port map( B1 => n57, B2 => n108, C1 => n59, C2 => n109, A 
                           => n110, ZN => n107);
   U185 : AOI22_X1 port map( A1 => REGISTERS_12_30_port, A2 => n62, B1 => 
                           REGISTERS_13_30_port, B2 => n63, ZN => n110);
   U186 : OAI221_X1 port map( B1 => n64, B2 => n111, C1 => n66, C2 => n112, A 
                           => n113, ZN => n106);
   U187 : AOI22_X1 port map( A1 => REGISTERS_8_30_port, A2 => n69, B1 => 
                           REGISTERS_9_30_port, B2 => n70, ZN => n113);
   U188 : OAI221_X1 port map( B1 => n71, B2 => n114, C1 => n73, C2 => n115, A 
                           => n116, ZN => n105);
   U189 : AOI22_X1 port map( A1 => REGISTERS_4_30_port, A2 => n76, B1 => 
                           REGISTERS_5_30_port, B2 => n77, ZN => n116);
   U190 : OAI221_X1 port map( B1 => n78, B2 => n117, C1 => n80, C2 => n118, A 
                           => n119, ZN => n104);
   U191 : AOI22_X1 port map( A1 => REGISTERS_0_30_port, A2 => n83, B1 => 
                           REGISTERS_1_30_port, B2 => n84, ZN => n119);
   U192 : NAND2_X1 port map( A1 => n120, A2 => n121, ZN => N2541);
   U193 : NOR4_X1 port map( A1 => n122, A2 => n123, A3 => n124, A4 => n125, ZN 
                           => n121);
   U194 : OAI221_X1 port map( B1 => n25, B2 => n126, C1 => n27, C2 => n127, A 
                           => n128, ZN => n125);
   U195 : AOI22_X1 port map( A1 => REGISTERS_28_29_port, A2 => n30, B1 => 
                           REGISTERS_29_29_port, B2 => n31, ZN => n128);
   U196 : OAI221_X1 port map( B1 => n32, B2 => n129, C1 => n34, C2 => n130, A 
                           => n131, ZN => n124);
   U197 : AOI22_X1 port map( A1 => REGISTERS_24_29_port, A2 => n37, B1 => 
                           REGISTERS_25_29_port, B2 => n38, ZN => n131);
   U198 : OAI221_X1 port map( B1 => n39, B2 => n132, C1 => n41, C2 => n133, A 
                           => n134, ZN => n123);
   U199 : AOI22_X1 port map( A1 => REGISTERS_20_29_port, A2 => n44, B1 => 
                           REGISTERS_21_29_port, B2 => n45, ZN => n134);
   U200 : OAI221_X1 port map( B1 => n46, B2 => n135, C1 => n48, C2 => n136, A 
                           => n137, ZN => n122);
   U201 : AOI22_X1 port map( A1 => REGISTERS_16_29_port, A2 => n51, B1 => 
                           REGISTERS_17_29_port, B2 => n52, ZN => n137);
   U202 : NOR4_X1 port map( A1 => n138, A2 => n139, A3 => n140, A4 => n141, ZN 
                           => n120);
   U203 : OAI221_X1 port map( B1 => n57, B2 => n142, C1 => n59, C2 => n143, A 
                           => n144, ZN => n141);
   U204 : AOI22_X1 port map( A1 => REGISTERS_12_29_port, A2 => n62, B1 => 
                           REGISTERS_13_29_port, B2 => n63, ZN => n144);
   U205 : OAI221_X1 port map( B1 => n64, B2 => n145, C1 => n66, C2 => n146, A 
                           => n147, ZN => n140);
   U206 : AOI22_X1 port map( A1 => REGISTERS_8_29_port, A2 => n69, B1 => 
                           REGISTERS_9_29_port, B2 => n70, ZN => n147);
   U207 : OAI221_X1 port map( B1 => n71, B2 => n148, C1 => n73, C2 => n149, A 
                           => n150, ZN => n139);
   U208 : AOI22_X1 port map( A1 => REGISTERS_4_29_port, A2 => n76, B1 => 
                           REGISTERS_5_29_port, B2 => n77, ZN => n150);
   U209 : OAI221_X1 port map( B1 => n78, B2 => n151, C1 => n80, C2 => n152, A 
                           => n153, ZN => n138);
   U210 : AOI22_X1 port map( A1 => REGISTERS_0_29_port, A2 => n83, B1 => 
                           REGISTERS_1_29_port, B2 => n84, ZN => n153);
   U211 : NAND2_X1 port map( A1 => n154, A2 => n155, ZN => N2539);
   U212 : NOR4_X1 port map( A1 => n156, A2 => n157, A3 => n158, A4 => n159, ZN 
                           => n155);
   U213 : OAI221_X1 port map( B1 => n25, B2 => n160, C1 => n27, C2 => n161, A 
                           => n162, ZN => n159);
   U214 : AOI22_X1 port map( A1 => REGISTERS_28_28_port, A2 => n30, B1 => 
                           REGISTERS_29_28_port, B2 => n31, ZN => n162);
   U215 : OAI221_X1 port map( B1 => n32, B2 => n163, C1 => n34, C2 => n164, A 
                           => n165, ZN => n158);
   U216 : AOI22_X1 port map( A1 => REGISTERS_24_28_port, A2 => n37, B1 => 
                           REGISTERS_25_28_port, B2 => n38, ZN => n165);
   U217 : OAI221_X1 port map( B1 => n39, B2 => n166, C1 => n41, C2 => n167, A 
                           => n168, ZN => n157);
   U218 : AOI22_X1 port map( A1 => REGISTERS_20_28_port, A2 => n44, B1 => 
                           REGISTERS_21_28_port, B2 => n45, ZN => n168);
   U219 : OAI221_X1 port map( B1 => n46, B2 => n169, C1 => n48, C2 => n170, A 
                           => n171, ZN => n156);
   U220 : AOI22_X1 port map( A1 => REGISTERS_16_28_port, A2 => n51, B1 => 
                           REGISTERS_17_28_port, B2 => n52, ZN => n171);
   U221 : NOR4_X1 port map( A1 => n172, A2 => n173, A3 => n174, A4 => n175, ZN 
                           => n154);
   U222 : OAI221_X1 port map( B1 => n57, B2 => n176, C1 => n59, C2 => n177, A 
                           => n178, ZN => n175);
   U223 : AOI22_X1 port map( A1 => REGISTERS_12_28_port, A2 => n62, B1 => 
                           REGISTERS_13_28_port, B2 => n63, ZN => n178);
   U224 : OAI221_X1 port map( B1 => n64, B2 => n179, C1 => n66, C2 => n180, A 
                           => n181, ZN => n174);
   U225 : AOI22_X1 port map( A1 => REGISTERS_8_28_port, A2 => n69, B1 => 
                           REGISTERS_9_28_port, B2 => n70, ZN => n181);
   U226 : OAI221_X1 port map( B1 => n71, B2 => n182, C1 => n73, C2 => n183, A 
                           => n184, ZN => n173);
   U227 : AOI22_X1 port map( A1 => REGISTERS_4_28_port, A2 => n76, B1 => 
                           REGISTERS_5_28_port, B2 => n77, ZN => n184);
   U228 : OAI221_X1 port map( B1 => n78, B2 => n185, C1 => n80, C2 => n186, A 
                           => n187, ZN => n172);
   U229 : AOI22_X1 port map( A1 => REGISTERS_0_28_port, A2 => n83, B1 => 
                           REGISTERS_1_28_port, B2 => n84, ZN => n187);
   U230 : NAND2_X1 port map( A1 => n188, A2 => n189, ZN => N2537);
   U231 : NOR4_X1 port map( A1 => n190, A2 => n191, A3 => n192, A4 => n193, ZN 
                           => n189);
   U232 : OAI221_X1 port map( B1 => n25, B2 => n194, C1 => n27, C2 => n195, A 
                           => n196, ZN => n193);
   U233 : AOI22_X1 port map( A1 => REGISTERS_28_27_port, A2 => n30, B1 => 
                           REGISTERS_29_27_port, B2 => n31, ZN => n196);
   U234 : OAI221_X1 port map( B1 => n32, B2 => n197, C1 => n34, C2 => n198, A 
                           => n199, ZN => n192);
   U235 : AOI22_X1 port map( A1 => REGISTERS_24_27_port, A2 => n37, B1 => 
                           REGISTERS_25_27_port, B2 => n38, ZN => n199);
   U236 : OAI221_X1 port map( B1 => n39, B2 => n200, C1 => n41, C2 => n201, A 
                           => n202, ZN => n191);
   U237 : AOI22_X1 port map( A1 => REGISTERS_20_27_port, A2 => n44, B1 => 
                           REGISTERS_21_27_port, B2 => n45, ZN => n202);
   U238 : OAI221_X1 port map( B1 => n46, B2 => n203, C1 => n48, C2 => n204, A 
                           => n205, ZN => n190);
   U239 : AOI22_X1 port map( A1 => REGISTERS_16_27_port, A2 => n51, B1 => 
                           REGISTERS_17_27_port, B2 => n52, ZN => n205);
   U240 : NOR4_X1 port map( A1 => n206, A2 => n207, A3 => n208, A4 => n209, ZN 
                           => n188);
   U241 : OAI221_X1 port map( B1 => n57, B2 => n210, C1 => n59, C2 => n211, A 
                           => n212, ZN => n209);
   U242 : AOI22_X1 port map( A1 => REGISTERS_12_27_port, A2 => n62, B1 => 
                           REGISTERS_13_27_port, B2 => n63, ZN => n212);
   U243 : OAI221_X1 port map( B1 => n64, B2 => n213, C1 => n66, C2 => n214, A 
                           => n215, ZN => n208);
   U244 : AOI22_X1 port map( A1 => REGISTERS_8_27_port, A2 => n69, B1 => 
                           REGISTERS_9_27_port, B2 => n70, ZN => n215);
   U245 : OAI221_X1 port map( B1 => n71, B2 => n216, C1 => n73, C2 => n217, A 
                           => n218, ZN => n207);
   U246 : AOI22_X1 port map( A1 => REGISTERS_4_27_port, A2 => n76, B1 => 
                           REGISTERS_5_27_port, B2 => n77, ZN => n218);
   U247 : OAI221_X1 port map( B1 => n78, B2 => n219, C1 => n80, C2 => n220, A 
                           => n221, ZN => n206);
   U248 : AOI22_X1 port map( A1 => REGISTERS_0_27_port, A2 => n83, B1 => 
                           REGISTERS_1_27_port, B2 => n84, ZN => n221);
   U249 : NAND2_X1 port map( A1 => n222, A2 => n223, ZN => N2535);
   U250 : NOR4_X1 port map( A1 => n224, A2 => n225, A3 => n226, A4 => n227, ZN 
                           => n223);
   U251 : OAI221_X1 port map( B1 => n25, B2 => n228, C1 => n27, C2 => n229, A 
                           => n230, ZN => n227);
   U252 : AOI22_X1 port map( A1 => REGISTERS_28_26_port, A2 => n30, B1 => 
                           REGISTERS_29_26_port, B2 => n31, ZN => n230);
   U253 : OAI221_X1 port map( B1 => n32, B2 => n231, C1 => n34, C2 => n232, A 
                           => n233, ZN => n226);
   U254 : AOI22_X1 port map( A1 => REGISTERS_24_26_port, A2 => n37, B1 => 
                           REGISTERS_25_26_port, B2 => n38, ZN => n233);
   U255 : OAI221_X1 port map( B1 => n39, B2 => n234, C1 => n41, C2 => n235, A 
                           => n236, ZN => n225);
   U256 : AOI22_X1 port map( A1 => REGISTERS_20_26_port, A2 => n44, B1 => 
                           REGISTERS_21_26_port, B2 => n45, ZN => n236);
   U257 : OAI221_X1 port map( B1 => n46, B2 => n237, C1 => n48, C2 => n238, A 
                           => n239, ZN => n224);
   U258 : AOI22_X1 port map( A1 => REGISTERS_16_26_port, A2 => n51, B1 => 
                           REGISTERS_17_26_port, B2 => n52, ZN => n239);
   U259 : NOR4_X1 port map( A1 => n240, A2 => n241, A3 => n242, A4 => n243, ZN 
                           => n222);
   U260 : OAI221_X1 port map( B1 => n57, B2 => n244, C1 => n59, C2 => n245, A 
                           => n246, ZN => n243);
   U261 : AOI22_X1 port map( A1 => REGISTERS_12_26_port, A2 => n62, B1 => 
                           REGISTERS_13_26_port, B2 => n63, ZN => n246);
   U262 : OAI221_X1 port map( B1 => n64, B2 => n247, C1 => n66, C2 => n248, A 
                           => n249, ZN => n242);
   U263 : AOI22_X1 port map( A1 => REGISTERS_8_26_port, A2 => n69, B1 => 
                           REGISTERS_9_26_port, B2 => n70, ZN => n249);
   U264 : OAI221_X1 port map( B1 => n71, B2 => n250, C1 => n73, C2 => n251, A 
                           => n252, ZN => n241);
   U265 : AOI22_X1 port map( A1 => REGISTERS_4_26_port, A2 => n76, B1 => 
                           REGISTERS_5_26_port, B2 => n77, ZN => n252);
   U266 : OAI221_X1 port map( B1 => n78, B2 => n253, C1 => n80, C2 => n254, A 
                           => n255, ZN => n240);
   U267 : AOI22_X1 port map( A1 => REGISTERS_0_26_port, A2 => n83, B1 => 
                           REGISTERS_1_26_port, B2 => n84, ZN => n255);
   U268 : NAND2_X1 port map( A1 => n256, A2 => n257, ZN => N2533);
   U269 : NOR4_X1 port map( A1 => n258, A2 => n259, A3 => n260, A4 => n261, ZN 
                           => n257);
   U270 : OAI221_X1 port map( B1 => n25, B2 => n262, C1 => n27, C2 => n263, A 
                           => n264, ZN => n261);
   U271 : AOI22_X1 port map( A1 => REGISTERS_28_25_port, A2 => n30, B1 => 
                           REGISTERS_29_25_port, B2 => n31, ZN => n264);
   U272 : OAI221_X1 port map( B1 => n32, B2 => n265, C1 => n34, C2 => n266, A 
                           => n267, ZN => n260);
   U273 : AOI22_X1 port map( A1 => REGISTERS_24_25_port, A2 => n37, B1 => 
                           REGISTERS_25_25_port, B2 => n38, ZN => n267);
   U274 : OAI221_X1 port map( B1 => n39, B2 => n268, C1 => n41, C2 => n269, A 
                           => n270, ZN => n259);
   U275 : AOI22_X1 port map( A1 => REGISTERS_20_25_port, A2 => n44, B1 => 
                           REGISTERS_21_25_port, B2 => n45, ZN => n270);
   U276 : OAI221_X1 port map( B1 => n46, B2 => n271, C1 => n48, C2 => n272, A 
                           => n273, ZN => n258);
   U277 : AOI22_X1 port map( A1 => REGISTERS_16_25_port, A2 => n51, B1 => 
                           REGISTERS_17_25_port, B2 => n52, ZN => n273);
   U278 : NOR4_X1 port map( A1 => n274, A2 => n275, A3 => n276, A4 => n277, ZN 
                           => n256);
   U279 : OAI221_X1 port map( B1 => n57, B2 => n278, C1 => n59, C2 => n279, A 
                           => n280, ZN => n277);
   U280 : AOI22_X1 port map( A1 => REGISTERS_12_25_port, A2 => n62, B1 => 
                           REGISTERS_13_25_port, B2 => n63, ZN => n280);
   U281 : OAI221_X1 port map( B1 => n64, B2 => n281, C1 => n66, C2 => n282, A 
                           => n283, ZN => n276);
   U282 : AOI22_X1 port map( A1 => REGISTERS_8_25_port, A2 => n69, B1 => 
                           REGISTERS_9_25_port, B2 => n70, ZN => n283);
   U283 : OAI221_X1 port map( B1 => n71, B2 => n284, C1 => n73, C2 => n285, A 
                           => n286, ZN => n275);
   U284 : AOI22_X1 port map( A1 => REGISTERS_4_25_port, A2 => n76, B1 => 
                           REGISTERS_5_25_port, B2 => n77, ZN => n286);
   U285 : OAI221_X1 port map( B1 => n78, B2 => n287, C1 => n80, C2 => n288, A 
                           => n289, ZN => n274);
   U286 : AOI22_X1 port map( A1 => REGISTERS_0_25_port, A2 => n83, B1 => 
                           REGISTERS_1_25_port, B2 => n84, ZN => n289);
   U287 : NAND2_X1 port map( A1 => n290, A2 => n291, ZN => N2531);
   U288 : NOR4_X1 port map( A1 => n292, A2 => n293, A3 => n294, A4 => n295, ZN 
                           => n291);
   U289 : OAI221_X1 port map( B1 => n25, B2 => n296, C1 => n27, C2 => n297, A 
                           => n298, ZN => n295);
   U290 : AOI22_X1 port map( A1 => REGISTERS_28_24_port, A2 => n30, B1 => 
                           REGISTERS_29_24_port, B2 => n31, ZN => n298);
   U291 : OAI221_X1 port map( B1 => n32, B2 => n299, C1 => n34, C2 => n300, A 
                           => n301, ZN => n294);
   U292 : AOI22_X1 port map( A1 => REGISTERS_24_24_port, A2 => n37, B1 => 
                           REGISTERS_25_24_port, B2 => n38, ZN => n301);
   U293 : OAI221_X1 port map( B1 => n39, B2 => n302, C1 => n41, C2 => n303, A 
                           => n304, ZN => n293);
   U294 : AOI22_X1 port map( A1 => REGISTERS_20_24_port, A2 => n44, B1 => 
                           REGISTERS_21_24_port, B2 => n45, ZN => n304);
   U295 : OAI221_X1 port map( B1 => n46, B2 => n305, C1 => n48, C2 => n306, A 
                           => n307, ZN => n292);
   U296 : AOI22_X1 port map( A1 => REGISTERS_16_24_port, A2 => n51, B1 => 
                           REGISTERS_17_24_port, B2 => n52, ZN => n307);
   U297 : NOR4_X1 port map( A1 => n308, A2 => n309, A3 => n310, A4 => n311, ZN 
                           => n290);
   U298 : OAI221_X1 port map( B1 => n57, B2 => n312, C1 => n59, C2 => n313, A 
                           => n314, ZN => n311);
   U299 : AOI22_X1 port map( A1 => REGISTERS_12_24_port, A2 => n62, B1 => 
                           REGISTERS_13_24_port, B2 => n63, ZN => n314);
   U300 : OAI221_X1 port map( B1 => n64, B2 => n315, C1 => n66, C2 => n316, A 
                           => n317, ZN => n310);
   U301 : AOI22_X1 port map( A1 => REGISTERS_8_24_port, A2 => n69, B1 => 
                           REGISTERS_9_24_port, B2 => n70, ZN => n317);
   U302 : OAI221_X1 port map( B1 => n71, B2 => n318, C1 => n73, C2 => n319, A 
                           => n320, ZN => n309);
   U303 : AOI22_X1 port map( A1 => REGISTERS_4_24_port, A2 => n76, B1 => 
                           REGISTERS_5_24_port, B2 => n77, ZN => n320);
   U304 : OAI221_X1 port map( B1 => n78, B2 => n321, C1 => n80, C2 => n322, A 
                           => n323, ZN => n308);
   U305 : AOI22_X1 port map( A1 => REGISTERS_0_24_port, A2 => n83, B1 => 
                           REGISTERS_1_24_port, B2 => n84, ZN => n323);
   U306 : NAND2_X1 port map( A1 => n324, A2 => n325, ZN => N2529);
   U307 : NOR4_X1 port map( A1 => n326, A2 => n327, A3 => n328, A4 => n329, ZN 
                           => n325);
   U308 : OAI221_X1 port map( B1 => n25, B2 => n330, C1 => n27, C2 => n331, A 
                           => n332, ZN => n329);
   U309 : AOI22_X1 port map( A1 => REGISTERS_28_23_port, A2 => n30, B1 => 
                           REGISTERS_29_23_port, B2 => n31, ZN => n332);
   U310 : OAI221_X1 port map( B1 => n32, B2 => n333, C1 => n34, C2 => n334, A 
                           => n335, ZN => n328);
   U311 : AOI22_X1 port map( A1 => REGISTERS_24_23_port, A2 => n37, B1 => 
                           REGISTERS_25_23_port, B2 => n38, ZN => n335);
   U312 : OAI221_X1 port map( B1 => n39, B2 => n336, C1 => n41, C2 => n337, A 
                           => n338, ZN => n327);
   U313 : AOI22_X1 port map( A1 => REGISTERS_20_23_port, A2 => n44, B1 => 
                           REGISTERS_21_23_port, B2 => n45, ZN => n338);
   U314 : OAI221_X1 port map( B1 => n46, B2 => n339, C1 => n48, C2 => n340, A 
                           => n341, ZN => n326);
   U315 : AOI22_X1 port map( A1 => REGISTERS_16_23_port, A2 => n51, B1 => 
                           REGISTERS_17_23_port, B2 => n52, ZN => n341);
   U316 : NOR4_X1 port map( A1 => n342, A2 => n343, A3 => n344, A4 => n345, ZN 
                           => n324);
   U317 : OAI221_X1 port map( B1 => n57, B2 => n346, C1 => n59, C2 => n347, A 
                           => n348, ZN => n345);
   U318 : AOI22_X1 port map( A1 => REGISTERS_12_23_port, A2 => n62, B1 => 
                           REGISTERS_13_23_port, B2 => n63, ZN => n348);
   U319 : OAI221_X1 port map( B1 => n64, B2 => n349, C1 => n66, C2 => n350, A 
                           => n351, ZN => n344);
   U320 : AOI22_X1 port map( A1 => REGISTERS_8_23_port, A2 => n69, B1 => 
                           REGISTERS_9_23_port, B2 => n70, ZN => n351);
   U321 : OAI221_X1 port map( B1 => n71, B2 => n352, C1 => n73, C2 => n353, A 
                           => n354, ZN => n343);
   U322 : AOI22_X1 port map( A1 => REGISTERS_4_23_port, A2 => n76, B1 => 
                           REGISTERS_5_23_port, B2 => n77, ZN => n354);
   U323 : OAI221_X1 port map( B1 => n78, B2 => n355, C1 => n80, C2 => n356, A 
                           => n357, ZN => n342);
   U324 : AOI22_X1 port map( A1 => REGISTERS_0_23_port, A2 => n83, B1 => 
                           REGISTERS_1_23_port, B2 => n84, ZN => n357);
   U325 : NAND2_X1 port map( A1 => n358, A2 => n359, ZN => N2527);
   U326 : NOR4_X1 port map( A1 => n360, A2 => n361, A3 => n362, A4 => n363, ZN 
                           => n359);
   U327 : OAI221_X1 port map( B1 => n25, B2 => n364, C1 => n27, C2 => n365, A 
                           => n366, ZN => n363);
   U328 : AOI22_X1 port map( A1 => REGISTERS_28_22_port, A2 => n30, B1 => 
                           REGISTERS_29_22_port, B2 => n31, ZN => n366);
   U329 : OAI221_X1 port map( B1 => n32, B2 => n367, C1 => n34, C2 => n368, A 
                           => n369, ZN => n362);
   U330 : AOI22_X1 port map( A1 => REGISTERS_24_22_port, A2 => n37, B1 => 
                           REGISTERS_25_22_port, B2 => n38, ZN => n369);
   U331 : OAI221_X1 port map( B1 => n39, B2 => n370, C1 => n41, C2 => n371, A 
                           => n372, ZN => n361);
   U332 : AOI22_X1 port map( A1 => REGISTERS_20_22_port, A2 => n44, B1 => 
                           REGISTERS_21_22_port, B2 => n45, ZN => n372);
   U333 : OAI221_X1 port map( B1 => n46, B2 => n373, C1 => n48, C2 => n374, A 
                           => n375, ZN => n360);
   U334 : AOI22_X1 port map( A1 => REGISTERS_16_22_port, A2 => n51, B1 => 
                           REGISTERS_17_22_port, B2 => n52, ZN => n375);
   U335 : NOR4_X1 port map( A1 => n376, A2 => n377, A3 => n378, A4 => n379, ZN 
                           => n358);
   U336 : OAI221_X1 port map( B1 => n57, B2 => n380, C1 => n59, C2 => n381, A 
                           => n382, ZN => n379);
   U337 : AOI22_X1 port map( A1 => REGISTERS_12_22_port, A2 => n62, B1 => 
                           REGISTERS_13_22_port, B2 => n63, ZN => n382);
   U338 : OAI221_X1 port map( B1 => n64, B2 => n383, C1 => n66, C2 => n384, A 
                           => n385, ZN => n378);
   U339 : AOI22_X1 port map( A1 => REGISTERS_8_22_port, A2 => n69, B1 => 
                           REGISTERS_9_22_port, B2 => n70, ZN => n385);
   U340 : OAI221_X1 port map( B1 => n71, B2 => n386, C1 => n73, C2 => n387, A 
                           => n388, ZN => n377);
   U341 : AOI22_X1 port map( A1 => REGISTERS_4_22_port, A2 => n76, B1 => 
                           REGISTERS_5_22_port, B2 => n77, ZN => n388);
   U342 : OAI221_X1 port map( B1 => n78, B2 => n389, C1 => n80, C2 => n390, A 
                           => n391, ZN => n376);
   U343 : AOI22_X1 port map( A1 => REGISTERS_0_22_port, A2 => n83, B1 => 
                           REGISTERS_1_22_port, B2 => n84, ZN => n391);
   U344 : NAND2_X1 port map( A1 => n392, A2 => n393, ZN => N2525);
   U345 : NOR4_X1 port map( A1 => n394, A2 => n395, A3 => n396, A4 => n397, ZN 
                           => n393);
   U346 : OAI221_X1 port map( B1 => n25, B2 => n398, C1 => n27, C2 => n399, A 
                           => n400, ZN => n397);
   U347 : AOI22_X1 port map( A1 => REGISTERS_28_21_port, A2 => n30, B1 => 
                           REGISTERS_29_21_port, B2 => n31, ZN => n400);
   U348 : OAI221_X1 port map( B1 => n32, B2 => n401, C1 => n34, C2 => n402, A 
                           => n403, ZN => n396);
   U349 : AOI22_X1 port map( A1 => REGISTERS_24_21_port, A2 => n37, B1 => 
                           REGISTERS_25_21_port, B2 => n38, ZN => n403);
   U350 : OAI221_X1 port map( B1 => n39, B2 => n404, C1 => n41, C2 => n405, A 
                           => n406, ZN => n395);
   U351 : AOI22_X1 port map( A1 => REGISTERS_20_21_port, A2 => n44, B1 => 
                           REGISTERS_21_21_port, B2 => n45, ZN => n406);
   U352 : OAI221_X1 port map( B1 => n46, B2 => n407, C1 => n48, C2 => n408, A 
                           => n409, ZN => n394);
   U353 : AOI22_X1 port map( A1 => REGISTERS_16_21_port, A2 => n51, B1 => 
                           REGISTERS_17_21_port, B2 => n52, ZN => n409);
   U354 : NOR4_X1 port map( A1 => n410, A2 => n411, A3 => n412, A4 => n413, ZN 
                           => n392);
   U355 : OAI221_X1 port map( B1 => n57, B2 => n414, C1 => n59, C2 => n415, A 
                           => n416, ZN => n413);
   U356 : AOI22_X1 port map( A1 => REGISTERS_12_21_port, A2 => n62, B1 => 
                           REGISTERS_13_21_port, B2 => n63, ZN => n416);
   U357 : OAI221_X1 port map( B1 => n64, B2 => n417, C1 => n66, C2 => n418, A 
                           => n419, ZN => n412);
   U358 : AOI22_X1 port map( A1 => REGISTERS_8_21_port, A2 => n69, B1 => 
                           REGISTERS_9_21_port, B2 => n70, ZN => n419);
   U359 : OAI221_X1 port map( B1 => n71, B2 => n420, C1 => n73, C2 => n421, A 
                           => n422, ZN => n411);
   U360 : AOI22_X1 port map( A1 => REGISTERS_4_21_port, A2 => n76, B1 => 
                           REGISTERS_5_21_port, B2 => n77, ZN => n422);
   U361 : OAI221_X1 port map( B1 => n78, B2 => n423, C1 => n80, C2 => n424, A 
                           => n425, ZN => n410);
   U362 : AOI22_X1 port map( A1 => REGISTERS_0_21_port, A2 => n83, B1 => 
                           REGISTERS_1_21_port, B2 => n84, ZN => n425);
   U363 : NAND2_X1 port map( A1 => n426, A2 => n427, ZN => N2523);
   U364 : NOR4_X1 port map( A1 => n428, A2 => n429, A3 => n430, A4 => n431, ZN 
                           => n427);
   U365 : OAI221_X1 port map( B1 => n25, B2 => n432, C1 => n27, C2 => n433, A 
                           => n434, ZN => n431);
   U366 : AOI22_X1 port map( A1 => REGISTERS_28_20_port, A2 => n30, B1 => 
                           REGISTERS_29_20_port, B2 => n31, ZN => n434);
   U367 : OAI221_X1 port map( B1 => n32, B2 => n435, C1 => n34, C2 => n436, A 
                           => n437, ZN => n430);
   U368 : AOI22_X1 port map( A1 => REGISTERS_24_20_port, A2 => n37, B1 => 
                           REGISTERS_25_20_port, B2 => n38, ZN => n437);
   U369 : OAI221_X1 port map( B1 => n39, B2 => n438, C1 => n41, C2 => n439, A 
                           => n440, ZN => n429);
   U370 : AOI22_X1 port map( A1 => REGISTERS_20_20_port, A2 => n44, B1 => 
                           REGISTERS_21_20_port, B2 => n45, ZN => n440);
   U371 : OAI221_X1 port map( B1 => n46, B2 => n441, C1 => n48, C2 => n442, A 
                           => n443, ZN => n428);
   U372 : AOI22_X1 port map( A1 => REGISTERS_16_20_port, A2 => n51, B1 => 
                           REGISTERS_17_20_port, B2 => n52, ZN => n443);
   U373 : NOR4_X1 port map( A1 => n444, A2 => n445, A3 => n446, A4 => n447, ZN 
                           => n426);
   U374 : OAI221_X1 port map( B1 => n57, B2 => n448, C1 => n59, C2 => n449, A 
                           => n450, ZN => n447);
   U375 : AOI22_X1 port map( A1 => REGISTERS_12_20_port, A2 => n62, B1 => 
                           REGISTERS_13_20_port, B2 => n63, ZN => n450);
   U376 : OAI221_X1 port map( B1 => n64, B2 => n451, C1 => n66, C2 => n452, A 
                           => n453, ZN => n446);
   U377 : AOI22_X1 port map( A1 => REGISTERS_8_20_port, A2 => n69, B1 => 
                           REGISTERS_9_20_port, B2 => n70, ZN => n453);
   U378 : OAI221_X1 port map( B1 => n71, B2 => n454, C1 => n73, C2 => n455, A 
                           => n456, ZN => n445);
   U379 : AOI22_X1 port map( A1 => REGISTERS_4_20_port, A2 => n76, B1 => 
                           REGISTERS_5_20_port, B2 => n77, ZN => n456);
   U380 : OAI221_X1 port map( B1 => n78, B2 => n457, C1 => n80, C2 => n458, A 
                           => n459, ZN => n444);
   U381 : AOI22_X1 port map( A1 => REGISTERS_0_20_port, A2 => n83, B1 => 
                           REGISTERS_1_20_port, B2 => n84, ZN => n459);
   U382 : NAND2_X1 port map( A1 => n460, A2 => n461, ZN => N2521);
   U383 : NOR4_X1 port map( A1 => n462, A2 => n463, A3 => n464, A4 => n465, ZN 
                           => n461);
   U384 : OAI221_X1 port map( B1 => n25, B2 => n466, C1 => n27, C2 => n467, A 
                           => n468, ZN => n465);
   U385 : AOI22_X1 port map( A1 => REGISTERS_28_19_port, A2 => n30, B1 => 
                           REGISTERS_29_19_port, B2 => n31, ZN => n468);
   U386 : OAI221_X1 port map( B1 => n32, B2 => n469, C1 => n34, C2 => n470, A 
                           => n471, ZN => n464);
   U387 : AOI22_X1 port map( A1 => REGISTERS_24_19_port, A2 => n37, B1 => 
                           REGISTERS_25_19_port, B2 => n38, ZN => n471);
   U388 : OAI221_X1 port map( B1 => n39, B2 => n472, C1 => n41, C2 => n473, A 
                           => n474, ZN => n463);
   U389 : AOI22_X1 port map( A1 => REGISTERS_20_19_port, A2 => n44, B1 => 
                           REGISTERS_21_19_port, B2 => n45, ZN => n474);
   U390 : OAI221_X1 port map( B1 => n46, B2 => n475, C1 => n48, C2 => n476, A 
                           => n477, ZN => n462);
   U391 : AOI22_X1 port map( A1 => REGISTERS_16_19_port, A2 => n51, B1 => 
                           REGISTERS_17_19_port, B2 => n52, ZN => n477);
   U392 : NOR4_X1 port map( A1 => n478, A2 => n479, A3 => n480, A4 => n481, ZN 
                           => n460);
   U393 : OAI221_X1 port map( B1 => n57, B2 => n482, C1 => n59, C2 => n483, A 
                           => n484, ZN => n481);
   U394 : AOI22_X1 port map( A1 => REGISTERS_12_19_port, A2 => n62, B1 => 
                           REGISTERS_13_19_port, B2 => n63, ZN => n484);
   U395 : OAI221_X1 port map( B1 => n64, B2 => n485, C1 => n66, C2 => n486, A 
                           => n487, ZN => n480);
   U396 : AOI22_X1 port map( A1 => REGISTERS_8_19_port, A2 => n69, B1 => 
                           REGISTERS_9_19_port, B2 => n70, ZN => n487);
   U397 : OAI221_X1 port map( B1 => n71, B2 => n488, C1 => n73, C2 => n489, A 
                           => n490, ZN => n479);
   U398 : AOI22_X1 port map( A1 => REGISTERS_4_19_port, A2 => n76, B1 => 
                           REGISTERS_5_19_port, B2 => n77, ZN => n490);
   U399 : OAI221_X1 port map( B1 => n78, B2 => n491, C1 => n80, C2 => n492, A 
                           => n493, ZN => n478);
   U400 : AOI22_X1 port map( A1 => REGISTERS_0_19_port, A2 => n83, B1 => 
                           REGISTERS_1_19_port, B2 => n84, ZN => n493);
   U401 : NAND2_X1 port map( A1 => n494, A2 => n495, ZN => N2519);
   U402 : NOR4_X1 port map( A1 => n496, A2 => n497, A3 => n498, A4 => n499, ZN 
                           => n495);
   U403 : OAI221_X1 port map( B1 => n25, B2 => n500, C1 => n27, C2 => n501, A 
                           => n502, ZN => n499);
   U404 : AOI22_X1 port map( A1 => REGISTERS_28_18_port, A2 => n30, B1 => 
                           REGISTERS_29_18_port, B2 => n31, ZN => n502);
   U405 : OAI221_X1 port map( B1 => n32, B2 => n503, C1 => n34, C2 => n504, A 
                           => n505, ZN => n498);
   U406 : AOI22_X1 port map( A1 => REGISTERS_24_18_port, A2 => n37, B1 => 
                           REGISTERS_25_18_port, B2 => n38, ZN => n505);
   U407 : OAI221_X1 port map( B1 => n39, B2 => n506, C1 => n41, C2 => n507, A 
                           => n508, ZN => n497);
   U408 : AOI22_X1 port map( A1 => REGISTERS_20_18_port, A2 => n44, B1 => 
                           REGISTERS_21_18_port, B2 => n45, ZN => n508);
   U409 : OAI221_X1 port map( B1 => n46, B2 => n509, C1 => n48, C2 => n510, A 
                           => n511, ZN => n496);
   U410 : AOI22_X1 port map( A1 => REGISTERS_16_18_port, A2 => n51, B1 => 
                           REGISTERS_17_18_port, B2 => n52, ZN => n511);
   U411 : NOR4_X1 port map( A1 => n512, A2 => n513, A3 => n514, A4 => n515, ZN 
                           => n494);
   U412 : OAI221_X1 port map( B1 => n57, B2 => n516, C1 => n59, C2 => n517, A 
                           => n518, ZN => n515);
   U413 : AOI22_X1 port map( A1 => REGISTERS_12_18_port, A2 => n62, B1 => 
                           REGISTERS_13_18_port, B2 => n63, ZN => n518);
   U414 : OAI221_X1 port map( B1 => n64, B2 => n519, C1 => n66, C2 => n520, A 
                           => n521, ZN => n514);
   U415 : AOI22_X1 port map( A1 => REGISTERS_8_18_port, A2 => n69, B1 => 
                           REGISTERS_9_18_port, B2 => n70, ZN => n521);
   U416 : OAI221_X1 port map( B1 => n71, B2 => n522, C1 => n73, C2 => n523, A 
                           => n524, ZN => n513);
   U417 : AOI22_X1 port map( A1 => REGISTERS_4_18_port, A2 => n76, B1 => 
                           REGISTERS_5_18_port, B2 => n77, ZN => n524);
   U418 : OAI221_X1 port map( B1 => n78, B2 => n525, C1 => n80, C2 => n526, A 
                           => n527, ZN => n512);
   U419 : AOI22_X1 port map( A1 => REGISTERS_0_18_port, A2 => n83, B1 => 
                           REGISTERS_1_18_port, B2 => n84, ZN => n527);
   U420 : NAND2_X1 port map( A1 => n528, A2 => n529, ZN => N2517);
   U421 : NOR4_X1 port map( A1 => n530, A2 => n531, A3 => n532, A4 => n533, ZN 
                           => n529);
   U422 : OAI221_X1 port map( B1 => n25, B2 => n534, C1 => n27, C2 => n535, A 
                           => n536, ZN => n533);
   U423 : AOI22_X1 port map( A1 => REGISTERS_28_17_port, A2 => n30, B1 => 
                           REGISTERS_29_17_port, B2 => n31, ZN => n536);
   U424 : OAI221_X1 port map( B1 => n32, B2 => n537, C1 => n34, C2 => n538, A 
                           => n539, ZN => n532);
   U425 : AOI22_X1 port map( A1 => REGISTERS_24_17_port, A2 => n37, B1 => 
                           REGISTERS_25_17_port, B2 => n38, ZN => n539);
   U426 : OAI221_X1 port map( B1 => n39, B2 => n540, C1 => n41, C2 => n541, A 
                           => n542, ZN => n531);
   U427 : AOI22_X1 port map( A1 => REGISTERS_20_17_port, A2 => n44, B1 => 
                           REGISTERS_21_17_port, B2 => n45, ZN => n542);
   U428 : OAI221_X1 port map( B1 => n46, B2 => n543, C1 => n48, C2 => n544, A 
                           => n545, ZN => n530);
   U429 : AOI22_X1 port map( A1 => REGISTERS_16_17_port, A2 => n51, B1 => 
                           REGISTERS_17_17_port, B2 => n52, ZN => n545);
   U430 : NOR4_X1 port map( A1 => n546, A2 => n547, A3 => n548, A4 => n549, ZN 
                           => n528);
   U431 : OAI221_X1 port map( B1 => n57, B2 => n550, C1 => n59, C2 => n551, A 
                           => n552, ZN => n549);
   U432 : AOI22_X1 port map( A1 => REGISTERS_12_17_port, A2 => n62, B1 => 
                           REGISTERS_13_17_port, B2 => n63, ZN => n552);
   U433 : OAI221_X1 port map( B1 => n64, B2 => n553, C1 => n66, C2 => n554, A 
                           => n555, ZN => n548);
   U434 : AOI22_X1 port map( A1 => REGISTERS_8_17_port, A2 => n69, B1 => 
                           REGISTERS_9_17_port, B2 => n70, ZN => n555);
   U435 : OAI221_X1 port map( B1 => n71, B2 => n556, C1 => n73, C2 => n557, A 
                           => n558, ZN => n547);
   U436 : AOI22_X1 port map( A1 => REGISTERS_4_17_port, A2 => n76, B1 => 
                           REGISTERS_5_17_port, B2 => n77, ZN => n558);
   U437 : OAI221_X1 port map( B1 => n78, B2 => n559, C1 => n80, C2 => n560, A 
                           => n561, ZN => n546);
   U438 : AOI22_X1 port map( A1 => REGISTERS_0_17_port, A2 => n83, B1 => 
                           REGISTERS_1_17_port, B2 => n84, ZN => n561);
   U439 : NAND2_X1 port map( A1 => n562, A2 => n563, ZN => N2515);
   U440 : NOR4_X1 port map( A1 => n564, A2 => n565, A3 => n566, A4 => n567, ZN 
                           => n563);
   U441 : OAI221_X1 port map( B1 => n25, B2 => n568, C1 => n27, C2 => n569, A 
                           => n570, ZN => n567);
   U442 : AOI22_X1 port map( A1 => REGISTERS_28_16_port, A2 => n30, B1 => 
                           REGISTERS_29_16_port, B2 => n31, ZN => n570);
   U443 : OAI221_X1 port map( B1 => n32, B2 => n571, C1 => n34, C2 => n572, A 
                           => n573, ZN => n566);
   U444 : AOI22_X1 port map( A1 => REGISTERS_24_16_port, A2 => n37, B1 => 
                           REGISTERS_25_16_port, B2 => n38, ZN => n573);
   U445 : OAI221_X1 port map( B1 => n39, B2 => n574, C1 => n41, C2 => n575, A 
                           => n576, ZN => n565);
   U446 : AOI22_X1 port map( A1 => REGISTERS_20_16_port, A2 => n44, B1 => 
                           REGISTERS_21_16_port, B2 => n45, ZN => n576);
   U447 : OAI221_X1 port map( B1 => n46, B2 => n577, C1 => n48, C2 => n578, A 
                           => n579, ZN => n564);
   U448 : AOI22_X1 port map( A1 => REGISTERS_16_16_port, A2 => n51, B1 => 
                           REGISTERS_17_16_port, B2 => n52, ZN => n579);
   U449 : NOR4_X1 port map( A1 => n580, A2 => n581, A3 => n582, A4 => n583, ZN 
                           => n562);
   U450 : OAI221_X1 port map( B1 => n57, B2 => n584, C1 => n59, C2 => n585, A 
                           => n586, ZN => n583);
   U451 : AOI22_X1 port map( A1 => REGISTERS_12_16_port, A2 => n62, B1 => 
                           REGISTERS_13_16_port, B2 => n63, ZN => n586);
   U452 : OAI221_X1 port map( B1 => n64, B2 => n587, C1 => n66, C2 => n588, A 
                           => n589, ZN => n582);
   U453 : AOI22_X1 port map( A1 => REGISTERS_8_16_port, A2 => n69, B1 => 
                           REGISTERS_9_16_port, B2 => n70, ZN => n589);
   U454 : OAI221_X1 port map( B1 => n71, B2 => n590, C1 => n73, C2 => n591, A 
                           => n592, ZN => n581);
   U455 : AOI22_X1 port map( A1 => REGISTERS_4_16_port, A2 => n76, B1 => 
                           REGISTERS_5_16_port, B2 => n77, ZN => n592);
   U456 : OAI221_X1 port map( B1 => n78, B2 => n593, C1 => n80, C2 => n594, A 
                           => n595, ZN => n580);
   U457 : AOI22_X1 port map( A1 => REGISTERS_0_16_port, A2 => n83, B1 => 
                           REGISTERS_1_16_port, B2 => n84, ZN => n595);
   U458 : NAND2_X1 port map( A1 => n596, A2 => n597, ZN => N2513);
   U459 : NOR4_X1 port map( A1 => n598, A2 => n599, A3 => n600, A4 => n601, ZN 
                           => n597);
   U460 : OAI221_X1 port map( B1 => n25, B2 => n602, C1 => n27, C2 => n603, A 
                           => n604, ZN => n601);
   U461 : AOI22_X1 port map( A1 => REGISTERS_28_15_port, A2 => n30, B1 => 
                           REGISTERS_29_15_port, B2 => n31, ZN => n604);
   U462 : OAI221_X1 port map( B1 => n32, B2 => n605, C1 => n34, C2 => n606, A 
                           => n607, ZN => n600);
   U463 : AOI22_X1 port map( A1 => REGISTERS_24_15_port, A2 => n37, B1 => 
                           REGISTERS_25_15_port, B2 => n38, ZN => n607);
   U464 : OAI221_X1 port map( B1 => n39, B2 => n608, C1 => n41, C2 => n609, A 
                           => n610, ZN => n599);
   U465 : AOI22_X1 port map( A1 => REGISTERS_20_15_port, A2 => n44, B1 => 
                           REGISTERS_21_15_port, B2 => n45, ZN => n610);
   U466 : OAI221_X1 port map( B1 => n46, B2 => n611, C1 => n48, C2 => n612, A 
                           => n613, ZN => n598);
   U467 : AOI22_X1 port map( A1 => REGISTERS_16_15_port, A2 => n51, B1 => 
                           REGISTERS_17_15_port, B2 => n52, ZN => n613);
   U468 : NOR4_X1 port map( A1 => n614, A2 => n615, A3 => n616, A4 => n617, ZN 
                           => n596);
   U469 : OAI221_X1 port map( B1 => n57, B2 => n618, C1 => n59, C2 => n619, A 
                           => n620, ZN => n617);
   U470 : AOI22_X1 port map( A1 => REGISTERS_12_15_port, A2 => n62, B1 => 
                           REGISTERS_13_15_port, B2 => n63, ZN => n620);
   U471 : OAI221_X1 port map( B1 => n64, B2 => n621, C1 => n66, C2 => n622, A 
                           => n623, ZN => n616);
   U472 : AOI22_X1 port map( A1 => REGISTERS_8_15_port, A2 => n69, B1 => 
                           REGISTERS_9_15_port, B2 => n70, ZN => n623);
   U473 : OAI221_X1 port map( B1 => n71, B2 => n624, C1 => n73, C2 => n625, A 
                           => n626, ZN => n615);
   U474 : AOI22_X1 port map( A1 => REGISTERS_4_15_port, A2 => n76, B1 => 
                           REGISTERS_5_15_port, B2 => n77, ZN => n626);
   U475 : OAI221_X1 port map( B1 => n78, B2 => n627, C1 => n80, C2 => n628, A 
                           => n629, ZN => n614);
   U476 : AOI22_X1 port map( A1 => REGISTERS_0_15_port, A2 => n83, B1 => 
                           REGISTERS_1_15_port, B2 => n84, ZN => n629);
   U477 : NAND2_X1 port map( A1 => n630, A2 => n631, ZN => N2511);
   U478 : NOR4_X1 port map( A1 => n632, A2 => n633, A3 => n634, A4 => n635, ZN 
                           => n631);
   U479 : OAI221_X1 port map( B1 => n25, B2 => n636, C1 => n27, C2 => n637, A 
                           => n638, ZN => n635);
   U480 : AOI22_X1 port map( A1 => REGISTERS_28_14_port, A2 => n30, B1 => 
                           REGISTERS_29_14_port, B2 => n31, ZN => n638);
   U481 : OAI221_X1 port map( B1 => n32, B2 => n639, C1 => n34, C2 => n640, A 
                           => n641, ZN => n634);
   U482 : AOI22_X1 port map( A1 => REGISTERS_24_14_port, A2 => n37, B1 => 
                           REGISTERS_25_14_port, B2 => n38, ZN => n641);
   U483 : OAI221_X1 port map( B1 => n39, B2 => n642, C1 => n41, C2 => n643, A 
                           => n644, ZN => n633);
   U484 : AOI22_X1 port map( A1 => REGISTERS_20_14_port, A2 => n44, B1 => 
                           REGISTERS_21_14_port, B2 => n45, ZN => n644);
   U485 : OAI221_X1 port map( B1 => n46, B2 => n645, C1 => n48, C2 => n646, A 
                           => n647, ZN => n632);
   U486 : AOI22_X1 port map( A1 => REGISTERS_16_14_port, A2 => n51, B1 => 
                           REGISTERS_17_14_port, B2 => n52, ZN => n647);
   U487 : NOR4_X1 port map( A1 => n648, A2 => n649, A3 => n650, A4 => n651, ZN 
                           => n630);
   U488 : OAI221_X1 port map( B1 => n57, B2 => n652, C1 => n59, C2 => n653, A 
                           => n654, ZN => n651);
   U489 : AOI22_X1 port map( A1 => REGISTERS_12_14_port, A2 => n62, B1 => 
                           REGISTERS_13_14_port, B2 => n63, ZN => n654);
   U490 : OAI221_X1 port map( B1 => n64, B2 => n655, C1 => n66, C2 => n656, A 
                           => n657, ZN => n650);
   U491 : AOI22_X1 port map( A1 => REGISTERS_8_14_port, A2 => n69, B1 => 
                           REGISTERS_9_14_port, B2 => n70, ZN => n657);
   U492 : OAI221_X1 port map( B1 => n71, B2 => n658, C1 => n73, C2 => n659, A 
                           => n660, ZN => n649);
   U493 : AOI22_X1 port map( A1 => REGISTERS_4_14_port, A2 => n76, B1 => 
                           REGISTERS_5_14_port, B2 => n77, ZN => n660);
   U494 : OAI221_X1 port map( B1 => n78, B2 => n661, C1 => n80, C2 => n662, A 
                           => n663, ZN => n648);
   U495 : AOI22_X1 port map( A1 => REGISTERS_0_14_port, A2 => n83, B1 => 
                           REGISTERS_1_14_port, B2 => n84, ZN => n663);
   U496 : NAND2_X1 port map( A1 => n664, A2 => n665, ZN => N2509);
   U497 : NOR4_X1 port map( A1 => n666, A2 => n667, A3 => n668, A4 => n669, ZN 
                           => n665);
   U498 : OAI221_X1 port map( B1 => n25, B2 => n670, C1 => n27, C2 => n671, A 
                           => n672, ZN => n669);
   U499 : AOI22_X1 port map( A1 => REGISTERS_28_13_port, A2 => n30, B1 => 
                           REGISTERS_29_13_port, B2 => n31, ZN => n672);
   U500 : OAI221_X1 port map( B1 => n32, B2 => n673, C1 => n34, C2 => n674, A 
                           => n675, ZN => n668);
   U501 : AOI22_X1 port map( A1 => REGISTERS_24_13_port, A2 => n37, B1 => 
                           REGISTERS_25_13_port, B2 => n38, ZN => n675);
   U502 : OAI221_X1 port map( B1 => n39, B2 => n676, C1 => n41, C2 => n677, A 
                           => n678, ZN => n667);
   U503 : AOI22_X1 port map( A1 => REGISTERS_20_13_port, A2 => n44, B1 => 
                           REGISTERS_21_13_port, B2 => n45, ZN => n678);
   U504 : OAI221_X1 port map( B1 => n46, B2 => n679, C1 => n48, C2 => n680, A 
                           => n681, ZN => n666);
   U505 : AOI22_X1 port map( A1 => REGISTERS_16_13_port, A2 => n51, B1 => 
                           REGISTERS_17_13_port, B2 => n52, ZN => n681);
   U506 : NOR4_X1 port map( A1 => n682, A2 => n683, A3 => n684, A4 => n685, ZN 
                           => n664);
   U507 : OAI221_X1 port map( B1 => n57, B2 => n686, C1 => n59, C2 => n687, A 
                           => n688, ZN => n685);
   U508 : AOI22_X1 port map( A1 => REGISTERS_12_13_port, A2 => n62, B1 => 
                           REGISTERS_13_13_port, B2 => n63, ZN => n688);
   U509 : OAI221_X1 port map( B1 => n64, B2 => n689, C1 => n66, C2 => n690, A 
                           => n691, ZN => n684);
   U510 : AOI22_X1 port map( A1 => REGISTERS_8_13_port, A2 => n69, B1 => 
                           REGISTERS_9_13_port, B2 => n70, ZN => n691);
   U511 : OAI221_X1 port map( B1 => n71, B2 => n692, C1 => n73, C2 => n693, A 
                           => n694, ZN => n683);
   U512 : AOI22_X1 port map( A1 => REGISTERS_4_13_port, A2 => n76, B1 => 
                           REGISTERS_5_13_port, B2 => n77, ZN => n694);
   U513 : OAI221_X1 port map( B1 => n78, B2 => n695, C1 => n80, C2 => n696, A 
                           => n697, ZN => n682);
   U514 : AOI22_X1 port map( A1 => REGISTERS_0_13_port, A2 => n83, B1 => 
                           REGISTERS_1_13_port, B2 => n84, ZN => n697);
   U515 : NAND2_X1 port map( A1 => n698, A2 => n699, ZN => N2507);
   U516 : NOR4_X1 port map( A1 => n700, A2 => n701, A3 => n702, A4 => n703, ZN 
                           => n699);
   U517 : OAI221_X1 port map( B1 => n25, B2 => n704, C1 => n27, C2 => n705, A 
                           => n706, ZN => n703);
   U518 : AOI22_X1 port map( A1 => REGISTERS_28_12_port, A2 => n30, B1 => 
                           REGISTERS_29_12_port, B2 => n31, ZN => n706);
   U519 : OAI221_X1 port map( B1 => n32, B2 => n707, C1 => n34, C2 => n708, A 
                           => n709, ZN => n702);
   U520 : AOI22_X1 port map( A1 => REGISTERS_24_12_port, A2 => n37, B1 => 
                           REGISTERS_25_12_port, B2 => n38, ZN => n709);
   U521 : OAI221_X1 port map( B1 => n39, B2 => n710, C1 => n41, C2 => n711, A 
                           => n712, ZN => n701);
   U522 : AOI22_X1 port map( A1 => REGISTERS_20_12_port, A2 => n44, B1 => 
                           REGISTERS_21_12_port, B2 => n45, ZN => n712);
   U523 : OAI221_X1 port map( B1 => n46, B2 => n713, C1 => n48, C2 => n714, A 
                           => n715, ZN => n700);
   U524 : AOI22_X1 port map( A1 => REGISTERS_16_12_port, A2 => n51, B1 => 
                           REGISTERS_17_12_port, B2 => n52, ZN => n715);
   U525 : NOR4_X1 port map( A1 => n716, A2 => n717, A3 => n718, A4 => n719, ZN 
                           => n698);
   U526 : OAI221_X1 port map( B1 => n57, B2 => n720, C1 => n59, C2 => n721, A 
                           => n722, ZN => n719);
   U527 : AOI22_X1 port map( A1 => REGISTERS_12_12_port, A2 => n62, B1 => 
                           REGISTERS_13_12_port, B2 => n63, ZN => n722);
   U528 : OAI221_X1 port map( B1 => n64, B2 => n723, C1 => n66, C2 => n724, A 
                           => n725, ZN => n718);
   U529 : AOI22_X1 port map( A1 => REGISTERS_8_12_port, A2 => n69, B1 => 
                           REGISTERS_9_12_port, B2 => n70, ZN => n725);
   U530 : OAI221_X1 port map( B1 => n71, B2 => n726, C1 => n73, C2 => n727, A 
                           => n728, ZN => n717);
   U531 : AOI22_X1 port map( A1 => REGISTERS_4_12_port, A2 => n76, B1 => 
                           REGISTERS_5_12_port, B2 => n77, ZN => n728);
   U532 : OAI221_X1 port map( B1 => n78, B2 => n729, C1 => n80, C2 => n730, A 
                           => n731, ZN => n716);
   U533 : AOI22_X1 port map( A1 => REGISTERS_0_12_port, A2 => n83, B1 => 
                           REGISTERS_1_12_port, B2 => n84, ZN => n731);
   U534 : NAND2_X1 port map( A1 => n732, A2 => n733, ZN => N2505);
   U535 : NOR4_X1 port map( A1 => n734, A2 => n735, A3 => n736, A4 => n737, ZN 
                           => n733);
   U536 : OAI221_X1 port map( B1 => n25, B2 => n738, C1 => n27, C2 => n739, A 
                           => n740, ZN => n737);
   U537 : AOI22_X1 port map( A1 => REGISTERS_28_11_port, A2 => n30, B1 => 
                           REGISTERS_29_11_port, B2 => n31, ZN => n740);
   U538 : OAI221_X1 port map( B1 => n32, B2 => n741, C1 => n34, C2 => n742, A 
                           => n743, ZN => n736);
   U539 : AOI22_X1 port map( A1 => REGISTERS_24_11_port, A2 => n37, B1 => 
                           REGISTERS_25_11_port, B2 => n38, ZN => n743);
   U540 : OAI221_X1 port map( B1 => n39, B2 => n744, C1 => n41, C2 => n745, A 
                           => n746, ZN => n735);
   U541 : AOI22_X1 port map( A1 => REGISTERS_20_11_port, A2 => n44, B1 => 
                           REGISTERS_21_11_port, B2 => n45, ZN => n746);
   U542 : OAI221_X1 port map( B1 => n46, B2 => n747, C1 => n48, C2 => n748, A 
                           => n749, ZN => n734);
   U543 : AOI22_X1 port map( A1 => REGISTERS_16_11_port, A2 => n51, B1 => 
                           REGISTERS_17_11_port, B2 => n52, ZN => n749);
   U544 : NOR4_X1 port map( A1 => n750, A2 => n751, A3 => n752, A4 => n753, ZN 
                           => n732);
   U545 : OAI221_X1 port map( B1 => n57, B2 => n754, C1 => n59, C2 => n755, A 
                           => n756, ZN => n753);
   U546 : AOI22_X1 port map( A1 => REGISTERS_12_11_port, A2 => n62, B1 => 
                           REGISTERS_13_11_port, B2 => n63, ZN => n756);
   U547 : OAI221_X1 port map( B1 => n64, B2 => n757, C1 => n66, C2 => n758, A 
                           => n759, ZN => n752);
   U548 : AOI22_X1 port map( A1 => REGISTERS_8_11_port, A2 => n69, B1 => 
                           REGISTERS_9_11_port, B2 => n70, ZN => n759);
   U549 : OAI221_X1 port map( B1 => n71, B2 => n760, C1 => n73, C2 => n761, A 
                           => n762, ZN => n751);
   U550 : AOI22_X1 port map( A1 => REGISTERS_4_11_port, A2 => n76, B1 => 
                           REGISTERS_5_11_port, B2 => n77, ZN => n762);
   U551 : OAI221_X1 port map( B1 => n78, B2 => n763, C1 => n80, C2 => n764, A 
                           => n765, ZN => n750);
   U552 : AOI22_X1 port map( A1 => REGISTERS_0_11_port, A2 => n83, B1 => 
                           REGISTERS_1_11_port, B2 => n84, ZN => n765);
   U553 : NAND2_X1 port map( A1 => n766, A2 => n767, ZN => N2503);
   U554 : NOR4_X1 port map( A1 => n768, A2 => n769, A3 => n770, A4 => n771, ZN 
                           => n767);
   U555 : OAI221_X1 port map( B1 => n25, B2 => n772, C1 => n27, C2 => n773, A 
                           => n774, ZN => n771);
   U556 : AOI22_X1 port map( A1 => REGISTERS_28_10_port, A2 => n30, B1 => 
                           REGISTERS_29_10_port, B2 => n31, ZN => n774);
   U557 : OAI221_X1 port map( B1 => n32, B2 => n775, C1 => n34, C2 => n776, A 
                           => n777, ZN => n770);
   U558 : AOI22_X1 port map( A1 => REGISTERS_24_10_port, A2 => n37, B1 => 
                           REGISTERS_25_10_port, B2 => n38, ZN => n777);
   U559 : OAI221_X1 port map( B1 => n39, B2 => n778, C1 => n41, C2 => n779, A 
                           => n780, ZN => n769);
   U560 : AOI22_X1 port map( A1 => REGISTERS_20_10_port, A2 => n44, B1 => 
                           REGISTERS_21_10_port, B2 => n45, ZN => n780);
   U561 : OAI221_X1 port map( B1 => n46, B2 => n781, C1 => n48, C2 => n782, A 
                           => n783, ZN => n768);
   U562 : AOI22_X1 port map( A1 => REGISTERS_16_10_port, A2 => n51, B1 => 
                           REGISTERS_17_10_port, B2 => n52, ZN => n783);
   U563 : NOR4_X1 port map( A1 => n784, A2 => n785, A3 => n786, A4 => n787, ZN 
                           => n766);
   U564 : OAI221_X1 port map( B1 => n57, B2 => n788, C1 => n59, C2 => n789, A 
                           => n790, ZN => n787);
   U565 : AOI22_X1 port map( A1 => REGISTERS_12_10_port, A2 => n62, B1 => 
                           REGISTERS_13_10_port, B2 => n63, ZN => n790);
   U566 : OAI221_X1 port map( B1 => n64, B2 => n791, C1 => n66, C2 => n792, A 
                           => n793, ZN => n786);
   U567 : AOI22_X1 port map( A1 => REGISTERS_8_10_port, A2 => n69, B1 => 
                           REGISTERS_9_10_port, B2 => n70, ZN => n793);
   U568 : OAI221_X1 port map( B1 => n71, B2 => n794, C1 => n73, C2 => n795, A 
                           => n796, ZN => n785);
   U569 : AOI22_X1 port map( A1 => REGISTERS_4_10_port, A2 => n76, B1 => 
                           REGISTERS_5_10_port, B2 => n77, ZN => n796);
   U570 : OAI221_X1 port map( B1 => n78, B2 => n797, C1 => n80, C2 => n798, A 
                           => n799, ZN => n784);
   U571 : AOI22_X1 port map( A1 => REGISTERS_0_10_port, A2 => n83, B1 => 
                           REGISTERS_1_10_port, B2 => n84, ZN => n799);
   U572 : NAND2_X1 port map( A1 => n800, A2 => n801, ZN => N2501);
   U573 : NOR4_X1 port map( A1 => n802, A2 => n803, A3 => n804, A4 => n805, ZN 
                           => n801);
   U574 : OAI221_X1 port map( B1 => n25, B2 => n806, C1 => n27, C2 => n807, A 
                           => n808, ZN => n805);
   U575 : AOI22_X1 port map( A1 => REGISTERS_28_9_port, A2 => n30, B1 => 
                           REGISTERS_29_9_port, B2 => n31, ZN => n808);
   U576 : OAI221_X1 port map( B1 => n32, B2 => n809, C1 => n34, C2 => n810, A 
                           => n811, ZN => n804);
   U577 : AOI22_X1 port map( A1 => REGISTERS_24_9_port, A2 => n37, B1 => 
                           REGISTERS_25_9_port, B2 => n38, ZN => n811);
   U578 : OAI221_X1 port map( B1 => n39, B2 => n812, C1 => n41, C2 => n813, A 
                           => n814, ZN => n803);
   U579 : AOI22_X1 port map( A1 => REGISTERS_20_9_port, A2 => n44, B1 => 
                           REGISTERS_21_9_port, B2 => n45, ZN => n814);
   U580 : OAI221_X1 port map( B1 => n46, B2 => n815, C1 => n48, C2 => n816, A 
                           => n817, ZN => n802);
   U581 : AOI22_X1 port map( A1 => REGISTERS_16_9_port, A2 => n51, B1 => 
                           REGISTERS_17_9_port, B2 => n52, ZN => n817);
   U582 : NOR4_X1 port map( A1 => n818, A2 => n819, A3 => n820, A4 => n821, ZN 
                           => n800);
   U583 : OAI221_X1 port map( B1 => n57, B2 => n822, C1 => n59, C2 => n823, A 
                           => n824, ZN => n821);
   U584 : AOI22_X1 port map( A1 => REGISTERS_12_9_port, A2 => n62, B1 => 
                           REGISTERS_13_9_port, B2 => n63, ZN => n824);
   U585 : OAI221_X1 port map( B1 => n64, B2 => n825, C1 => n66, C2 => n826, A 
                           => n827, ZN => n820);
   U586 : AOI22_X1 port map( A1 => REGISTERS_8_9_port, A2 => n69, B1 => 
                           REGISTERS_9_9_port, B2 => n70, ZN => n827);
   U587 : OAI221_X1 port map( B1 => n71, B2 => n828, C1 => n73, C2 => n829, A 
                           => n830, ZN => n819);
   U588 : AOI22_X1 port map( A1 => REGISTERS_4_9_port, A2 => n76, B1 => 
                           REGISTERS_5_9_port, B2 => n77, ZN => n830);
   U589 : OAI221_X1 port map( B1 => n78, B2 => n831, C1 => n80, C2 => n832, A 
                           => n833, ZN => n818);
   U590 : AOI22_X1 port map( A1 => REGISTERS_0_9_port, A2 => n83, B1 => 
                           REGISTERS_1_9_port, B2 => n84, ZN => n833);
   U591 : NAND2_X1 port map( A1 => n834, A2 => n835, ZN => N2499);
   U592 : NOR4_X1 port map( A1 => n836, A2 => n837, A3 => n838, A4 => n839, ZN 
                           => n835);
   U593 : OAI221_X1 port map( B1 => n25, B2 => n840, C1 => n27, C2 => n841, A 
                           => n842, ZN => n839);
   U594 : AOI22_X1 port map( A1 => REGISTERS_28_8_port, A2 => n30, B1 => 
                           REGISTERS_29_8_port, B2 => n31, ZN => n842);
   U595 : OAI221_X1 port map( B1 => n32, B2 => n843, C1 => n34, C2 => n844, A 
                           => n845, ZN => n838);
   U596 : AOI22_X1 port map( A1 => REGISTERS_24_8_port, A2 => n37, B1 => 
                           REGISTERS_25_8_port, B2 => n38, ZN => n845);
   U597 : OAI221_X1 port map( B1 => n39, B2 => n846, C1 => n41, C2 => n847, A 
                           => n848, ZN => n837);
   U598 : AOI22_X1 port map( A1 => REGISTERS_20_8_port, A2 => n44, B1 => 
                           REGISTERS_21_8_port, B2 => n45, ZN => n848);
   U599 : OAI221_X1 port map( B1 => n46, B2 => n849, C1 => n48, C2 => n850, A 
                           => n851, ZN => n836);
   U600 : AOI22_X1 port map( A1 => REGISTERS_16_8_port, A2 => n51, B1 => 
                           REGISTERS_17_8_port, B2 => n52, ZN => n851);
   U601 : NOR4_X1 port map( A1 => n852, A2 => n853, A3 => n854, A4 => n855, ZN 
                           => n834);
   U602 : OAI221_X1 port map( B1 => n57, B2 => n856, C1 => n59, C2 => n857, A 
                           => n858, ZN => n855);
   U603 : AOI22_X1 port map( A1 => REGISTERS_12_8_port, A2 => n62, B1 => 
                           REGISTERS_13_8_port, B2 => n63, ZN => n858);
   U604 : OAI221_X1 port map( B1 => n64, B2 => n859, C1 => n66, C2 => n860, A 
                           => n861, ZN => n854);
   U605 : AOI22_X1 port map( A1 => REGISTERS_8_8_port, A2 => n69, B1 => 
                           REGISTERS_9_8_port, B2 => n70, ZN => n861);
   U606 : OAI221_X1 port map( B1 => n71, B2 => n862, C1 => n73, C2 => n863, A 
                           => n864, ZN => n853);
   U607 : AOI22_X1 port map( A1 => REGISTERS_4_8_port, A2 => n76, B1 => 
                           REGISTERS_5_8_port, B2 => n77, ZN => n864);
   U608 : OAI221_X1 port map( B1 => n78, B2 => n865, C1 => n80, C2 => n866, A 
                           => n867, ZN => n852);
   U609 : AOI22_X1 port map( A1 => REGISTERS_0_8_port, A2 => n83, B1 => 
                           REGISTERS_1_8_port, B2 => n84, ZN => n867);
   U610 : NAND2_X1 port map( A1 => n868, A2 => n869, ZN => N2497);
   U611 : NOR4_X1 port map( A1 => n870, A2 => n871, A3 => n872, A4 => n873, ZN 
                           => n869);
   U612 : OAI221_X1 port map( B1 => n25, B2 => n874, C1 => n27, C2 => n875, A 
                           => n876, ZN => n873);
   U613 : AOI22_X1 port map( A1 => REGISTERS_28_7_port, A2 => n30, B1 => 
                           REGISTERS_29_7_port, B2 => n31, ZN => n876);
   U614 : OAI221_X1 port map( B1 => n32, B2 => n877, C1 => n34, C2 => n878, A 
                           => n879, ZN => n872);
   U615 : AOI22_X1 port map( A1 => REGISTERS_24_7_port, A2 => n37, B1 => 
                           REGISTERS_25_7_port, B2 => n38, ZN => n879);
   U616 : OAI221_X1 port map( B1 => n39, B2 => n880, C1 => n41, C2 => n881, A 
                           => n882, ZN => n871);
   U617 : AOI22_X1 port map( A1 => REGISTERS_20_7_port, A2 => n44, B1 => 
                           REGISTERS_21_7_port, B2 => n45, ZN => n882);
   U618 : OAI221_X1 port map( B1 => n46, B2 => n883, C1 => n48, C2 => n884, A 
                           => n885, ZN => n870);
   U619 : AOI22_X1 port map( A1 => REGISTERS_16_7_port, A2 => n51, B1 => 
                           REGISTERS_17_7_port, B2 => n52, ZN => n885);
   U620 : NOR4_X1 port map( A1 => n886, A2 => n887, A3 => n888, A4 => n889, ZN 
                           => n868);
   U621 : OAI221_X1 port map( B1 => n57, B2 => n890, C1 => n59, C2 => n891, A 
                           => n892, ZN => n889);
   U622 : AOI22_X1 port map( A1 => REGISTERS_12_7_port, A2 => n62, B1 => 
                           REGISTERS_13_7_port, B2 => n63, ZN => n892);
   U623 : OAI221_X1 port map( B1 => n64, B2 => n893, C1 => n66, C2 => n894, A 
                           => n895, ZN => n888);
   U624 : AOI22_X1 port map( A1 => REGISTERS_8_7_port, A2 => n69, B1 => 
                           REGISTERS_9_7_port, B2 => n70, ZN => n895);
   U625 : OAI221_X1 port map( B1 => n71, B2 => n896, C1 => n73, C2 => n897, A 
                           => n898, ZN => n887);
   U626 : AOI22_X1 port map( A1 => REGISTERS_4_7_port, A2 => n76, B1 => 
                           REGISTERS_5_7_port, B2 => n77, ZN => n898);
   U627 : OAI221_X1 port map( B1 => n78, B2 => n899, C1 => n80, C2 => n900, A 
                           => n901, ZN => n886);
   U628 : AOI22_X1 port map( A1 => REGISTERS_0_7_port, A2 => n83, B1 => 
                           REGISTERS_1_7_port, B2 => n84, ZN => n901);
   U629 : NAND2_X1 port map( A1 => n902, A2 => n903, ZN => N2495);
   U630 : NOR4_X1 port map( A1 => n904, A2 => n905, A3 => n906, A4 => n907, ZN 
                           => n903);
   U631 : OAI221_X1 port map( B1 => n25, B2 => n908, C1 => n27, C2 => n909, A 
                           => n910, ZN => n907);
   U632 : AOI22_X1 port map( A1 => REGISTERS_28_6_port, A2 => n30, B1 => 
                           REGISTERS_29_6_port, B2 => n31, ZN => n910);
   U633 : OAI221_X1 port map( B1 => n32, B2 => n911, C1 => n34, C2 => n912, A 
                           => n913, ZN => n906);
   U634 : AOI22_X1 port map( A1 => REGISTERS_24_6_port, A2 => n37, B1 => 
                           REGISTERS_25_6_port, B2 => n38, ZN => n913);
   U635 : OAI221_X1 port map( B1 => n39, B2 => n914, C1 => n41, C2 => n915, A 
                           => n916, ZN => n905);
   U636 : AOI22_X1 port map( A1 => REGISTERS_20_6_port, A2 => n44, B1 => 
                           REGISTERS_21_6_port, B2 => n45, ZN => n916);
   U637 : OAI221_X1 port map( B1 => n46, B2 => n917, C1 => n48, C2 => n918, A 
                           => n919, ZN => n904);
   U638 : AOI22_X1 port map( A1 => REGISTERS_16_6_port, A2 => n51, B1 => 
                           REGISTERS_17_6_port, B2 => n52, ZN => n919);
   U639 : NOR4_X1 port map( A1 => n920, A2 => n921, A3 => n922, A4 => n923, ZN 
                           => n902);
   U640 : OAI221_X1 port map( B1 => n57, B2 => n924, C1 => n59, C2 => n925, A 
                           => n926, ZN => n923);
   U641 : AOI22_X1 port map( A1 => REGISTERS_12_6_port, A2 => n62, B1 => 
                           REGISTERS_13_6_port, B2 => n63, ZN => n926);
   U642 : OAI221_X1 port map( B1 => n64, B2 => n927, C1 => n66, C2 => n928, A 
                           => n929, ZN => n922);
   U643 : AOI22_X1 port map( A1 => REGISTERS_8_6_port, A2 => n69, B1 => 
                           REGISTERS_9_6_port, B2 => n70, ZN => n929);
   U644 : OAI221_X1 port map( B1 => n71, B2 => n930, C1 => n73, C2 => n931, A 
                           => n932, ZN => n921);
   U645 : AOI22_X1 port map( A1 => REGISTERS_4_6_port, A2 => n76, B1 => 
                           REGISTERS_5_6_port, B2 => n77, ZN => n932);
   U646 : OAI221_X1 port map( B1 => n78, B2 => n933, C1 => n80, C2 => n934, A 
                           => n935, ZN => n920);
   U647 : AOI22_X1 port map( A1 => REGISTERS_0_6_port, A2 => n83, B1 => 
                           REGISTERS_1_6_port, B2 => n84, ZN => n935);
   U648 : NAND2_X1 port map( A1 => n936, A2 => n937, ZN => N2493);
   U649 : NOR4_X1 port map( A1 => n938, A2 => n939, A3 => n940, A4 => n941, ZN 
                           => n937);
   U650 : OAI221_X1 port map( B1 => n25, B2 => n942, C1 => n27, C2 => n943, A 
                           => n944, ZN => n941);
   U651 : AOI22_X1 port map( A1 => REGISTERS_28_5_port, A2 => n30, B1 => 
                           REGISTERS_29_5_port, B2 => n31, ZN => n944);
   U652 : OAI221_X1 port map( B1 => n32, B2 => n945, C1 => n34, C2 => n946, A 
                           => n947, ZN => n940);
   U653 : AOI22_X1 port map( A1 => REGISTERS_24_5_port, A2 => n37, B1 => 
                           REGISTERS_25_5_port, B2 => n38, ZN => n947);
   U654 : OAI221_X1 port map( B1 => n39, B2 => n948, C1 => n41, C2 => n949, A 
                           => n950, ZN => n939);
   U655 : AOI22_X1 port map( A1 => REGISTERS_20_5_port, A2 => n44, B1 => 
                           REGISTERS_21_5_port, B2 => n45, ZN => n950);
   U656 : OAI221_X1 port map( B1 => n46, B2 => n951, C1 => n48, C2 => n952, A 
                           => n953, ZN => n938);
   U657 : AOI22_X1 port map( A1 => REGISTERS_16_5_port, A2 => n51, B1 => 
                           REGISTERS_17_5_port, B2 => n52, ZN => n953);
   U658 : NOR4_X1 port map( A1 => n954, A2 => n955, A3 => n956, A4 => n957, ZN 
                           => n936);
   U659 : OAI221_X1 port map( B1 => n57, B2 => n958, C1 => n59, C2 => n959, A 
                           => n960, ZN => n957);
   U660 : AOI22_X1 port map( A1 => REGISTERS_12_5_port, A2 => n62, B1 => 
                           REGISTERS_13_5_port, B2 => n63, ZN => n960);
   U661 : OAI221_X1 port map( B1 => n64, B2 => n961, C1 => n66, C2 => n962, A 
                           => n963, ZN => n956);
   U662 : AOI22_X1 port map( A1 => REGISTERS_8_5_port, A2 => n69, B1 => 
                           REGISTERS_9_5_port, B2 => n70, ZN => n963);
   U663 : OAI221_X1 port map( B1 => n71, B2 => n964, C1 => n73, C2 => n965, A 
                           => n966, ZN => n955);
   U664 : AOI22_X1 port map( A1 => REGISTERS_4_5_port, A2 => n76, B1 => 
                           REGISTERS_5_5_port, B2 => n77, ZN => n966);
   U665 : OAI221_X1 port map( B1 => n78, B2 => n967, C1 => n80, C2 => n968, A 
                           => n969, ZN => n954);
   U666 : AOI22_X1 port map( A1 => REGISTERS_0_5_port, A2 => n83, B1 => 
                           REGISTERS_1_5_port, B2 => n84, ZN => n969);
   U667 : NAND2_X1 port map( A1 => n970, A2 => n971, ZN => N2491);
   U668 : NOR4_X1 port map( A1 => n972, A2 => n973, A3 => n974, A4 => n975, ZN 
                           => n971);
   U669 : OAI221_X1 port map( B1 => n25, B2 => n976, C1 => n27, C2 => n977, A 
                           => n978, ZN => n975);
   U670 : AOI22_X1 port map( A1 => REGISTERS_28_4_port, A2 => n30, B1 => 
                           REGISTERS_29_4_port, B2 => n31, ZN => n978);
   U671 : OAI221_X1 port map( B1 => n32, B2 => n979, C1 => n34, C2 => n980, A 
                           => n981, ZN => n974);
   U672 : AOI22_X1 port map( A1 => REGISTERS_24_4_port, A2 => n37, B1 => 
                           REGISTERS_25_4_port, B2 => n38, ZN => n981);
   U673 : OAI221_X1 port map( B1 => n39, B2 => n982, C1 => n41, C2 => n983, A 
                           => n984, ZN => n973);
   U674 : AOI22_X1 port map( A1 => REGISTERS_20_4_port, A2 => n44, B1 => 
                           REGISTERS_21_4_port, B2 => n45, ZN => n984);
   U675 : OAI221_X1 port map( B1 => n46, B2 => n985, C1 => n48, C2 => n986, A 
                           => n987, ZN => n972);
   U676 : AOI22_X1 port map( A1 => REGISTERS_16_4_port, A2 => n51, B1 => 
                           REGISTERS_17_4_port, B2 => n52, ZN => n987);
   U677 : NOR4_X1 port map( A1 => n988, A2 => n989, A3 => n990, A4 => n991, ZN 
                           => n970);
   U678 : OAI221_X1 port map( B1 => n57, B2 => n992, C1 => n59, C2 => n993, A 
                           => n994, ZN => n991);
   U679 : AOI22_X1 port map( A1 => REGISTERS_12_4_port, A2 => n62, B1 => 
                           REGISTERS_13_4_port, B2 => n63, ZN => n994);
   U680 : OAI221_X1 port map( B1 => n64, B2 => n995, C1 => n66, C2 => n996, A 
                           => n997, ZN => n990);
   U681 : AOI22_X1 port map( A1 => REGISTERS_8_4_port, A2 => n69, B1 => 
                           REGISTERS_9_4_port, B2 => n70, ZN => n997);
   U682 : OAI221_X1 port map( B1 => n71, B2 => n998, C1 => n73, C2 => n999, A 
                           => n1000, ZN => n989);
   U683 : AOI22_X1 port map( A1 => REGISTERS_4_4_port, A2 => n76, B1 => 
                           REGISTERS_5_4_port, B2 => n77, ZN => n1000);
   U684 : OAI221_X1 port map( B1 => n78, B2 => n1001, C1 => n80, C2 => n1002, A
                           => n1003, ZN => n988);
   U685 : AOI22_X1 port map( A1 => REGISTERS_0_4_port, A2 => n83, B1 => 
                           REGISTERS_1_4_port, B2 => n84, ZN => n1003);
   U686 : NAND2_X1 port map( A1 => n1004, A2 => n1005, ZN => N2489);
   U687 : NOR4_X1 port map( A1 => n1006, A2 => n1007, A3 => n1008, A4 => n1009,
                           ZN => n1005);
   U688 : OAI221_X1 port map( B1 => n25, B2 => n1010, C1 => n27, C2 => n1011, A
                           => n1012, ZN => n1009);
   U689 : AOI22_X1 port map( A1 => REGISTERS_28_3_port, A2 => n30, B1 => 
                           REGISTERS_29_3_port, B2 => n31, ZN => n1012);
   U690 : OAI221_X1 port map( B1 => n32, B2 => n1013, C1 => n34, C2 => n1014, A
                           => n1015, ZN => n1008);
   U691 : AOI22_X1 port map( A1 => REGISTERS_24_3_port, A2 => n37, B1 => 
                           REGISTERS_25_3_port, B2 => n38, ZN => n1015);
   U692 : OAI221_X1 port map( B1 => n39, B2 => n1016, C1 => n41, C2 => n1017, A
                           => n1018, ZN => n1007);
   U693 : AOI22_X1 port map( A1 => REGISTERS_20_3_port, A2 => n44, B1 => 
                           REGISTERS_21_3_port, B2 => n45, ZN => n1018);
   U694 : OAI221_X1 port map( B1 => n46, B2 => n1019, C1 => n48, C2 => n1020, A
                           => n1021, ZN => n1006);
   U695 : AOI22_X1 port map( A1 => REGISTERS_16_3_port, A2 => n51, B1 => 
                           REGISTERS_17_3_port, B2 => n52, ZN => n1021);
   U696 : NOR4_X1 port map( A1 => n1022, A2 => n1023, A3 => n1024, A4 => n1025,
                           ZN => n1004);
   U697 : OAI221_X1 port map( B1 => n57, B2 => n1026, C1 => n59, C2 => n1027, A
                           => n1028, ZN => n1025);
   U698 : AOI22_X1 port map( A1 => REGISTERS_12_3_port, A2 => n62, B1 => 
                           REGISTERS_13_3_port, B2 => n63, ZN => n1028);
   U699 : OAI221_X1 port map( B1 => n64, B2 => n1029, C1 => n66, C2 => n1030, A
                           => n1031, ZN => n1024);
   U700 : AOI22_X1 port map( A1 => REGISTERS_8_3_port, A2 => n69, B1 => 
                           REGISTERS_9_3_port, B2 => n70, ZN => n1031);
   U701 : OAI221_X1 port map( B1 => n71, B2 => n1032, C1 => n73, C2 => n1033, A
                           => n1034, ZN => n1023);
   U702 : AOI22_X1 port map( A1 => REGISTERS_4_3_port, A2 => n76, B1 => 
                           REGISTERS_5_3_port, B2 => n77, ZN => n1034);
   U703 : OAI221_X1 port map( B1 => n78, B2 => n1035, C1 => n80, C2 => n1036, A
                           => n1037, ZN => n1022);
   U704 : AOI22_X1 port map( A1 => REGISTERS_0_3_port, A2 => n83, B1 => 
                           REGISTERS_1_3_port, B2 => n84, ZN => n1037);
   U705 : NAND2_X1 port map( A1 => n1038, A2 => n1039, ZN => N2487);
   U706 : NOR4_X1 port map( A1 => n1040, A2 => n1041, A3 => n1042, A4 => n1043,
                           ZN => n1039);
   U707 : OAI221_X1 port map( B1 => n25, B2 => n1044, C1 => n27, C2 => n1045, A
                           => n1046, ZN => n1043);
   U708 : AOI22_X1 port map( A1 => REGISTERS_28_2_port, A2 => n30, B1 => 
                           REGISTERS_29_2_port, B2 => n31, ZN => n1046);
   U709 : OAI221_X1 port map( B1 => n32, B2 => n1047, C1 => n34, C2 => n1048, A
                           => n1049, ZN => n1042);
   U710 : AOI22_X1 port map( A1 => REGISTERS_24_2_port, A2 => n37, B1 => 
                           REGISTERS_25_2_port, B2 => n38, ZN => n1049);
   U711 : OAI221_X1 port map( B1 => n39, B2 => n1050, C1 => n41, C2 => n1051, A
                           => n1052, ZN => n1041);
   U712 : AOI22_X1 port map( A1 => REGISTERS_20_2_port, A2 => n44, B1 => 
                           REGISTERS_21_2_port, B2 => n45, ZN => n1052);
   U713 : OAI221_X1 port map( B1 => n46, B2 => n1053, C1 => n48, C2 => n1054, A
                           => n1055, ZN => n1040);
   U714 : AOI22_X1 port map( A1 => REGISTERS_16_2_port, A2 => n51, B1 => 
                           REGISTERS_17_2_port, B2 => n52, ZN => n1055);
   U715 : NOR4_X1 port map( A1 => n1056, A2 => n1057, A3 => n1058, A4 => n1059,
                           ZN => n1038);
   U716 : OAI221_X1 port map( B1 => n57, B2 => n1060, C1 => n59, C2 => n1061, A
                           => n1062, ZN => n1059);
   U717 : AOI22_X1 port map( A1 => REGISTERS_12_2_port, A2 => n62, B1 => 
                           REGISTERS_13_2_port, B2 => n63, ZN => n1062);
   U718 : OAI221_X1 port map( B1 => n64, B2 => n1063, C1 => n66, C2 => n1064, A
                           => n1065, ZN => n1058);
   U719 : AOI22_X1 port map( A1 => REGISTERS_8_2_port, A2 => n69, B1 => 
                           REGISTERS_9_2_port, B2 => n70, ZN => n1065);
   U720 : OAI221_X1 port map( B1 => n71, B2 => n1066, C1 => n73, C2 => n1067, A
                           => n1068, ZN => n1057);
   U721 : AOI22_X1 port map( A1 => REGISTERS_4_2_port, A2 => n76, B1 => 
                           REGISTERS_5_2_port, B2 => n77, ZN => n1068);
   U722 : OAI221_X1 port map( B1 => n78, B2 => n1069, C1 => n80, C2 => n1070, A
                           => n1071, ZN => n1056);
   U723 : AOI22_X1 port map( A1 => REGISTERS_0_2_port, A2 => n83, B1 => 
                           REGISTERS_1_2_port, B2 => n84, ZN => n1071);
   U724 : NAND2_X1 port map( A1 => n1072, A2 => n1073, ZN => N2485);
   U725 : NOR4_X1 port map( A1 => n1074, A2 => n1075, A3 => n1076, A4 => n1077,
                           ZN => n1073);
   U726 : OAI221_X1 port map( B1 => n25, B2 => n1078, C1 => n27, C2 => n1079, A
                           => n1080, ZN => n1077);
   U727 : AOI22_X1 port map( A1 => REGISTERS_28_1_port, A2 => n30, B1 => 
                           REGISTERS_29_1_port, B2 => n31, ZN => n1080);
   U728 : OAI221_X1 port map( B1 => n32, B2 => n1081, C1 => n34, C2 => n1082, A
                           => n1083, ZN => n1076);
   U729 : AOI22_X1 port map( A1 => REGISTERS_24_1_port, A2 => n37, B1 => 
                           REGISTERS_25_1_port, B2 => n38, ZN => n1083);
   U730 : OAI221_X1 port map( B1 => n39, B2 => n1084, C1 => n41, C2 => n1085, A
                           => n1086, ZN => n1075);
   U731 : AOI22_X1 port map( A1 => REGISTERS_20_1_port, A2 => n44, B1 => 
                           REGISTERS_21_1_port, B2 => n45, ZN => n1086);
   U732 : OAI221_X1 port map( B1 => n46, B2 => n1087, C1 => n48, C2 => n1088, A
                           => n1089, ZN => n1074);
   U733 : AOI22_X1 port map( A1 => REGISTERS_16_1_port, A2 => n51, B1 => 
                           REGISTERS_17_1_port, B2 => n52, ZN => n1089);
   U734 : NOR4_X1 port map( A1 => n1090, A2 => n1091, A3 => n1092, A4 => n1093,
                           ZN => n1072);
   U735 : OAI221_X1 port map( B1 => n57, B2 => n1094, C1 => n59, C2 => n1095, A
                           => n1096, ZN => n1093);
   U736 : AOI22_X1 port map( A1 => REGISTERS_12_1_port, A2 => n62, B1 => 
                           REGISTERS_13_1_port, B2 => n63, ZN => n1096);
   U737 : OAI221_X1 port map( B1 => n64, B2 => n1097, C1 => n66, C2 => n1098, A
                           => n1099, ZN => n1092);
   U738 : AOI22_X1 port map( A1 => REGISTERS_8_1_port, A2 => n69, B1 => 
                           REGISTERS_9_1_port, B2 => n70, ZN => n1099);
   U739 : OAI221_X1 port map( B1 => n71, B2 => n1100, C1 => n73, C2 => n1101, A
                           => n1102, ZN => n1091);
   U740 : AOI22_X1 port map( A1 => REGISTERS_4_1_port, A2 => n76, B1 => 
                           REGISTERS_5_1_port, B2 => n77, ZN => n1102);
   U741 : OAI221_X1 port map( B1 => n78, B2 => n1103, C1 => n80, C2 => n1104, A
                           => n1105, ZN => n1090);
   U742 : AOI22_X1 port map( A1 => REGISTERS_0_1_port, A2 => n83, B1 => 
                           REGISTERS_1_1_port, B2 => n84, ZN => n1105);
   U743 : NAND2_X1 port map( A1 => n1106, A2 => n1107, ZN => N2483);
   U744 : NOR4_X1 port map( A1 => n1108, A2 => n1109, A3 => n1110, A4 => n1111,
                           ZN => n1107);
   U745 : OAI221_X1 port map( B1 => n25, B2 => n1112, C1 => n27, C2 => n1113, A
                           => n1114, ZN => n1111);
   U746 : AOI22_X1 port map( A1 => REGISTERS_28_0_port, A2 => n30, B1 => 
                           REGISTERS_29_0_port, B2 => n31, ZN => n1114);
   U747 : OAI221_X1 port map( B1 => n32, B2 => n1119, C1 => n34, C2 => n1120, A
                           => n1121, ZN => n1110);
   U748 : AOI22_X1 port map( A1 => REGISTERS_24_0_port, A2 => n37, B1 => 
                           REGISTERS_25_0_port, B2 => n38, ZN => n1121);
   U749 : AND3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(3), ZN => n1115);
   U750 : AND3_X1 port map( A1 => ADD_RD2(4), A2 => n1124, A3 => ADD_RD2(3), ZN
                           => n1117);
   U751 : OAI221_X1 port map( B1 => n39, B2 => n1125, C1 => n41, C2 => n1126, A
                           => n1127, ZN => n1109);
   U752 : AOI22_X1 port map( A1 => REGISTERS_20_0_port, A2 => n44, B1 => 
                           REGISTERS_21_0_port, B2 => n45, ZN => n1127);
   U753 : OAI221_X1 port map( B1 => n46, B2 => n1130, C1 => n48, C2 => n1131, A
                           => n1132, ZN => n1108);
   U754 : AOI22_X1 port map( A1 => REGISTERS_16_0_port, A2 => n51, B1 => 
                           REGISTERS_17_0_port, B2 => n52, ZN => n1132);
   U755 : AND3_X1 port map( A1 => ADD_RD2(4), A2 => n1133, A3 => ADD_RD2(0), ZN
                           => n1128);
   U756 : AND3_X1 port map( A1 => n1124, A2 => n1133, A3 => ADD_RD2(4), ZN => 
                           n1129);
   U757 : NOR4_X1 port map( A1 => n1134, A2 => n1135, A3 => n1136, A4 => n1137,
                           ZN => n1106);
   U758 : OAI221_X1 port map( B1 => n57, B2 => n1138, C1 => n59, C2 => n1139, A
                           => n1140, ZN => n1137);
   U759 : AOI22_X1 port map( A1 => REGISTERS_12_0_port, A2 => n62, B1 => 
                           REGISTERS_13_0_port, B2 => n63, ZN => n1140);
   U760 : OAI221_X1 port map( B1 => n64, B2 => n1143, C1 => n66, C2 => n1144, A
                           => n1145, ZN => n1136);
   U761 : AOI22_X1 port map( A1 => REGISTERS_8_0_port, A2 => n69, B1 => 
                           REGISTERS_9_0_port, B2 => n70, ZN => n1145);
   U762 : NOR3_X1 port map( A1 => n1124, A2 => ADD_RD2(4), A3 => n1133, ZN => 
                           n1141);
   U763 : NOR3_X1 port map( A1 => ADD_RD2(0), A2 => ADD_RD2(4), A3 => n1133, ZN
                           => n1142);
   U764 : INV_X1 port map( A => ADD_RD2(3), ZN => n1133);
   U765 : OAI221_X1 port map( B1 => n71, B2 => n1146, C1 => n73, C2 => n1147, A
                           => n1148, ZN => n1135);
   U766 : AOI22_X1 port map( A1 => REGISTERS_4_0_port, A2 => n76, B1 => 
                           REGISTERS_5_0_port, B2 => n77, ZN => n1148);
   U767 : AND3_X1 port map( A1 => n1151, A2 => n1152, A3 => ADD_RD2(2), ZN => 
                           n1116);
   U768 : AND3_X1 port map( A1 => ADD_RD2(1), A2 => n1151, A3 => ADD_RD2(2), ZN
                           => n1118);
   U769 : OAI221_X1 port map( B1 => n78, B2 => n1153, C1 => n80, C2 => n1154, A
                           => n1155, ZN => n1134);
   U770 : AOI22_X1 port map( A1 => REGISTERS_0_0_port, A2 => n83, B1 => 
                           REGISTERS_1_0_port, B2 => n84, ZN => n1155);
   U771 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => n1124, ZN
                           => n1149);
   U772 : INV_X1 port map( A => ADD_RD2(0), ZN => n1124);
   U773 : INV_X1 port map( A => ADD_RD2(1), ZN => n1152);
   U774 : NOR3_X1 port map( A1 => ADD_RD2(3), A2 => ADD_RD2(4), A3 => 
                           ADD_RD2(0), ZN => n1150);
   U775 : NAND2_X1 port map( A1 => n1156, A2 => n1157, ZN => N2481);
   U776 : NOR4_X1 port map( A1 => n1158, A2 => n1159, A3 => n1160, A4 => n1161,
                           ZN => n1157);
   U777 : OAI221_X1 port map( B1 => n26, B2 => n1162, C1 => n28, C2 => n1163, A
                           => n1164, ZN => n1161);
   U778 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_31_port, B1 => 
                           n1166, B2 => REGISTERS_29_31_port, ZN => n1164);
   U779 : INV_X1 port map( A => REGISTERS_31_31_port, ZN => n28);
   U780 : INV_X1 port map( A => REGISTERS_30_31_port, ZN => n26);
   U781 : OAI221_X1 port map( B1 => n33, B2 => n1167, C1 => n35, C2 => n1168, A
                           => n1169, ZN => n1160);
   U782 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_31_port, B1 => 
                           n1171, B2 => REGISTERS_25_31_port, ZN => n1169);
   U783 : INV_X1 port map( A => REGISTERS_27_31_port, ZN => n35);
   U784 : INV_X1 port map( A => REGISTERS_26_31_port, ZN => n33);
   U785 : OAI221_X1 port map( B1 => n40, B2 => n1172, C1 => n42, C2 => n1173, A
                           => n1174, ZN => n1159);
   U786 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_31_port, B1 => 
                           n1176, B2 => REGISTERS_21_31_port, ZN => n1174);
   U787 : INV_X1 port map( A => REGISTERS_23_31_port, ZN => n42);
   U788 : INV_X1 port map( A => REGISTERS_22_31_port, ZN => n40);
   U789 : OAI221_X1 port map( B1 => n47, B2 => n1177, C1 => n49, C2 => n1178, A
                           => n1179, ZN => n1158);
   U790 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_31_port, B1 => 
                           n1181, B2 => REGISTERS_17_31_port, ZN => n1179);
   U791 : INV_X1 port map( A => REGISTERS_19_31_port, ZN => n49);
   U792 : INV_X1 port map( A => REGISTERS_18_31_port, ZN => n47);
   U793 : NOR4_X1 port map( A1 => n1182, A2 => n1183, A3 => n1184, A4 => n1185,
                           ZN => n1156);
   U794 : OAI221_X1 port map( B1 => n58, B2 => n1186, C1 => n60, C2 => n1187, A
                           => n1188, ZN => n1185);
   U795 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_31_port, B1 => 
                           n1190, B2 => REGISTERS_13_31_port, ZN => n1188);
   U796 : INV_X1 port map( A => REGISTERS_15_31_port, ZN => n60);
   U797 : INV_X1 port map( A => REGISTERS_14_31_port, ZN => n58);
   U798 : OAI221_X1 port map( B1 => n65, B2 => n1191, C1 => n67, C2 => n1192, A
                           => n1193, ZN => n1184);
   U799 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_31_port, B1 => 
                           n1195, B2 => REGISTERS_9_31_port, ZN => n1193);
   U800 : INV_X1 port map( A => REGISTERS_11_31_port, ZN => n67);
   U801 : INV_X1 port map( A => REGISTERS_10_31_port, ZN => n65);
   U802 : OAI221_X1 port map( B1 => n72, B2 => n1196, C1 => n74, C2 => n1197, A
                           => n1198, ZN => n1183);
   U803 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_31_port, B1 => 
                           n1200, B2 => REGISTERS_5_31_port, ZN => n1198);
   U804 : INV_X1 port map( A => REGISTERS_7_31_port, ZN => n74);
   U805 : INV_X1 port map( A => REGISTERS_6_31_port, ZN => n72);
   U806 : OAI221_X1 port map( B1 => n79, B2 => n1201, C1 => n81, C2 => n1202, A
                           => n1203, ZN => n1182);
   U807 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_31_port, B1 => 
                           n1205, B2 => REGISTERS_1_31_port, ZN => n1203);
   U808 : INV_X1 port map( A => REGISTERS_3_31_port, ZN => n81);
   U809 : INV_X1 port map( A => REGISTERS_2_31_port, ZN => n79);
   U810 : OR2_X1 port map( A1 => RD1, A2 => n85, ZN => N2480);
   U811 : NAND2_X1 port map( A1 => n1206, A2 => n1207, ZN => N2479);
   U812 : NOR4_X1 port map( A1 => n1208, A2 => n1209, A3 => n1210, A4 => n1211,
                           ZN => n1207);
   U813 : OAI221_X1 port map( B1 => n92, B2 => n1162, C1 => n93, C2 => n1163, A
                           => n1212, ZN => n1211);
   U814 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_30_port, B1 => 
                           n1166, B2 => REGISTERS_29_30_port, ZN => n1212);
   U815 : INV_X1 port map( A => REGISTERS_31_30_port, ZN => n93);
   U816 : INV_X1 port map( A => REGISTERS_30_30_port, ZN => n92);
   U817 : OAI221_X1 port map( B1 => n95, B2 => n1167, C1 => n96, C2 => n1168, A
                           => n1213, ZN => n1210);
   U818 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_30_port, B1 => 
                           n1171, B2 => REGISTERS_25_30_port, ZN => n1213);
   U819 : INV_X1 port map( A => REGISTERS_27_30_port, ZN => n96);
   U820 : INV_X1 port map( A => REGISTERS_26_30_port, ZN => n95);
   U821 : OAI221_X1 port map( B1 => n98, B2 => n1172, C1 => n99, C2 => n1173, A
                           => n1214, ZN => n1209);
   U822 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_30_port, B1 => 
                           n1176, B2 => REGISTERS_21_30_port, ZN => n1214);
   U823 : INV_X1 port map( A => REGISTERS_23_30_port, ZN => n99);
   U824 : INV_X1 port map( A => REGISTERS_22_30_port, ZN => n98);
   U825 : OAI221_X1 port map( B1 => n101, B2 => n1177, C1 => n102, C2 => n1178,
                           A => n1215, ZN => n1208);
   U826 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_30_port, B1 => 
                           n1181, B2 => REGISTERS_17_30_port, ZN => n1215);
   U827 : INV_X1 port map( A => REGISTERS_19_30_port, ZN => n102);
   U828 : INV_X1 port map( A => REGISTERS_18_30_port, ZN => n101);
   U829 : NOR4_X1 port map( A1 => n1216, A2 => n1217, A3 => n1218, A4 => n1219,
                           ZN => n1206);
   U830 : OAI221_X1 port map( B1 => n108, B2 => n1186, C1 => n109, C2 => n1187,
                           A => n1220, ZN => n1219);
   U831 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_30_port, B1 => 
                           n1190, B2 => REGISTERS_13_30_port, ZN => n1220);
   U832 : INV_X1 port map( A => REGISTERS_15_30_port, ZN => n109);
   U833 : INV_X1 port map( A => REGISTERS_14_30_port, ZN => n108);
   U834 : OAI221_X1 port map( B1 => n111, B2 => n1191, C1 => n112, C2 => n1192,
                           A => n1221, ZN => n1218);
   U835 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_30_port, B1 => 
                           n1195, B2 => REGISTERS_9_30_port, ZN => n1221);
   U836 : INV_X1 port map( A => REGISTERS_11_30_port, ZN => n112);
   U837 : INV_X1 port map( A => REGISTERS_10_30_port, ZN => n111);
   U838 : OAI221_X1 port map( B1 => n114, B2 => n1196, C1 => n115, C2 => n1197,
                           A => n1222, ZN => n1217);
   U839 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_30_port, B1 => 
                           n1200, B2 => REGISTERS_5_30_port, ZN => n1222);
   U840 : INV_X1 port map( A => REGISTERS_7_30_port, ZN => n115);
   U841 : INV_X1 port map( A => REGISTERS_6_30_port, ZN => n114);
   U842 : OAI221_X1 port map( B1 => n117, B2 => n1201, C1 => n118, C2 => n1202,
                           A => n1223, ZN => n1216);
   U843 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_30_port, B1 => 
                           n1205, B2 => REGISTERS_1_30_port, ZN => n1223);
   U844 : INV_X1 port map( A => REGISTERS_3_30_port, ZN => n118);
   U845 : INV_X1 port map( A => REGISTERS_2_30_port, ZN => n117);
   U846 : NAND2_X1 port map( A1 => n1224, A2 => n1225, ZN => N2477);
   U847 : NOR4_X1 port map( A1 => n1226, A2 => n1227, A3 => n1228, A4 => n1229,
                           ZN => n1225);
   U848 : OAI221_X1 port map( B1 => n126, B2 => n1162, C1 => n127, C2 => n1163,
                           A => n1230, ZN => n1229);
   U849 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_29_port, B1 => 
                           n1166, B2 => REGISTERS_29_29_port, ZN => n1230);
   U850 : INV_X1 port map( A => REGISTERS_31_29_port, ZN => n127);
   U851 : INV_X1 port map( A => REGISTERS_30_29_port, ZN => n126);
   U852 : OAI221_X1 port map( B1 => n129, B2 => n1167, C1 => n130, C2 => n1168,
                           A => n1231, ZN => n1228);
   U853 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_29_port, B1 => 
                           n1171, B2 => REGISTERS_25_29_port, ZN => n1231);
   U854 : INV_X1 port map( A => REGISTERS_27_29_port, ZN => n130);
   U855 : INV_X1 port map( A => REGISTERS_26_29_port, ZN => n129);
   U856 : OAI221_X1 port map( B1 => n132, B2 => n1172, C1 => n133, C2 => n1173,
                           A => n1232, ZN => n1227);
   U857 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_29_port, B1 => 
                           n1176, B2 => REGISTERS_21_29_port, ZN => n1232);
   U858 : INV_X1 port map( A => REGISTERS_23_29_port, ZN => n133);
   U859 : INV_X1 port map( A => REGISTERS_22_29_port, ZN => n132);
   U860 : OAI221_X1 port map( B1 => n135, B2 => n1177, C1 => n136, C2 => n1178,
                           A => n1233, ZN => n1226);
   U861 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_29_port, B1 => 
                           n1181, B2 => REGISTERS_17_29_port, ZN => n1233);
   U862 : INV_X1 port map( A => REGISTERS_19_29_port, ZN => n136);
   U863 : INV_X1 port map( A => REGISTERS_18_29_port, ZN => n135);
   U864 : NOR4_X1 port map( A1 => n1234, A2 => n1235, A3 => n1236, A4 => n1237,
                           ZN => n1224);
   U865 : OAI221_X1 port map( B1 => n142, B2 => n1186, C1 => n143, C2 => n1187,
                           A => n1238, ZN => n1237);
   U866 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_29_port, B1 => 
                           n1190, B2 => REGISTERS_13_29_port, ZN => n1238);
   U867 : INV_X1 port map( A => REGISTERS_15_29_port, ZN => n143);
   U868 : INV_X1 port map( A => REGISTERS_14_29_port, ZN => n142);
   U869 : OAI221_X1 port map( B1 => n145, B2 => n1191, C1 => n146, C2 => n1192,
                           A => n1239, ZN => n1236);
   U870 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_29_port, B1 => 
                           n1195, B2 => REGISTERS_9_29_port, ZN => n1239);
   U871 : INV_X1 port map( A => REGISTERS_11_29_port, ZN => n146);
   U872 : INV_X1 port map( A => REGISTERS_10_29_port, ZN => n145);
   U873 : OAI221_X1 port map( B1 => n148, B2 => n1196, C1 => n149, C2 => n1197,
                           A => n1240, ZN => n1235);
   U874 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_29_port, B1 => 
                           n1200, B2 => REGISTERS_5_29_port, ZN => n1240);
   U875 : INV_X1 port map( A => REGISTERS_7_29_port, ZN => n149);
   U876 : INV_X1 port map( A => REGISTERS_6_29_port, ZN => n148);
   U877 : OAI221_X1 port map( B1 => n151, B2 => n1201, C1 => n152, C2 => n1202,
                           A => n1241, ZN => n1234);
   U878 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_29_port, B1 => 
                           n1205, B2 => REGISTERS_1_29_port, ZN => n1241);
   U879 : INV_X1 port map( A => REGISTERS_3_29_port, ZN => n152);
   U880 : INV_X1 port map( A => REGISTERS_2_29_port, ZN => n151);
   U881 : NAND2_X1 port map( A1 => n1242, A2 => n1243, ZN => N2475);
   U882 : NOR4_X1 port map( A1 => n1244, A2 => n1245, A3 => n1246, A4 => n1247,
                           ZN => n1243);
   U883 : OAI221_X1 port map( B1 => n160, B2 => n1162, C1 => n161, C2 => n1163,
                           A => n1248, ZN => n1247);
   U884 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_28_port, B1 => 
                           n1166, B2 => REGISTERS_29_28_port, ZN => n1248);
   U885 : INV_X1 port map( A => REGISTERS_31_28_port, ZN => n161);
   U886 : INV_X1 port map( A => REGISTERS_30_28_port, ZN => n160);
   U887 : OAI221_X1 port map( B1 => n163, B2 => n1167, C1 => n164, C2 => n1168,
                           A => n1249, ZN => n1246);
   U888 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_28_port, B1 => 
                           n1171, B2 => REGISTERS_25_28_port, ZN => n1249);
   U889 : INV_X1 port map( A => REGISTERS_27_28_port, ZN => n164);
   U890 : INV_X1 port map( A => REGISTERS_26_28_port, ZN => n163);
   U891 : OAI221_X1 port map( B1 => n166, B2 => n1172, C1 => n167, C2 => n1173,
                           A => n1250, ZN => n1245);
   U892 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_28_port, B1 => 
                           n1176, B2 => REGISTERS_21_28_port, ZN => n1250);
   U893 : INV_X1 port map( A => REGISTERS_23_28_port, ZN => n167);
   U894 : INV_X1 port map( A => REGISTERS_22_28_port, ZN => n166);
   U895 : OAI221_X1 port map( B1 => n169, B2 => n1177, C1 => n170, C2 => n1178,
                           A => n1251, ZN => n1244);
   U896 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_28_port, B1 => 
                           n1181, B2 => REGISTERS_17_28_port, ZN => n1251);
   U897 : INV_X1 port map( A => REGISTERS_19_28_port, ZN => n170);
   U898 : INV_X1 port map( A => REGISTERS_18_28_port, ZN => n169);
   U899 : NOR4_X1 port map( A1 => n1252, A2 => n1253, A3 => n1254, A4 => n1255,
                           ZN => n1242);
   U900 : OAI221_X1 port map( B1 => n176, B2 => n1186, C1 => n177, C2 => n1187,
                           A => n1256, ZN => n1255);
   U901 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_28_port, B1 => 
                           n1190, B2 => REGISTERS_13_28_port, ZN => n1256);
   U902 : INV_X1 port map( A => REGISTERS_15_28_port, ZN => n177);
   U903 : INV_X1 port map( A => REGISTERS_14_28_port, ZN => n176);
   U904 : OAI221_X1 port map( B1 => n179, B2 => n1191, C1 => n180, C2 => n1192,
                           A => n1257, ZN => n1254);
   U905 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_28_port, B1 => 
                           n1195, B2 => REGISTERS_9_28_port, ZN => n1257);
   U906 : INV_X1 port map( A => REGISTERS_11_28_port, ZN => n180);
   U907 : INV_X1 port map( A => REGISTERS_10_28_port, ZN => n179);
   U908 : OAI221_X1 port map( B1 => n182, B2 => n1196, C1 => n183, C2 => n1197,
                           A => n1258, ZN => n1253);
   U909 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_28_port, B1 => 
                           n1200, B2 => REGISTERS_5_28_port, ZN => n1258);
   U910 : INV_X1 port map( A => REGISTERS_7_28_port, ZN => n183);
   U911 : INV_X1 port map( A => REGISTERS_6_28_port, ZN => n182);
   U912 : OAI221_X1 port map( B1 => n185, B2 => n1201, C1 => n186, C2 => n1202,
                           A => n1259, ZN => n1252);
   U913 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_28_port, B1 => 
                           n1205, B2 => REGISTERS_1_28_port, ZN => n1259);
   U914 : INV_X1 port map( A => REGISTERS_3_28_port, ZN => n186);
   U915 : INV_X1 port map( A => REGISTERS_2_28_port, ZN => n185);
   U916 : NAND2_X1 port map( A1 => n1260, A2 => n1261, ZN => N2473);
   U917 : NOR4_X1 port map( A1 => n1262, A2 => n1263, A3 => n1264, A4 => n1265,
                           ZN => n1261);
   U918 : OAI221_X1 port map( B1 => n194, B2 => n1162, C1 => n195, C2 => n1163,
                           A => n1266, ZN => n1265);
   U919 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_27_port, B1 => 
                           n1166, B2 => REGISTERS_29_27_port, ZN => n1266);
   U920 : INV_X1 port map( A => REGISTERS_31_27_port, ZN => n195);
   U921 : INV_X1 port map( A => REGISTERS_30_27_port, ZN => n194);
   U922 : OAI221_X1 port map( B1 => n197, B2 => n1167, C1 => n198, C2 => n1168,
                           A => n1267, ZN => n1264);
   U923 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_27_port, B1 => 
                           n1171, B2 => REGISTERS_25_27_port, ZN => n1267);
   U924 : INV_X1 port map( A => REGISTERS_27_27_port, ZN => n198);
   U925 : INV_X1 port map( A => REGISTERS_26_27_port, ZN => n197);
   U926 : OAI221_X1 port map( B1 => n200, B2 => n1172, C1 => n201, C2 => n1173,
                           A => n1268, ZN => n1263);
   U927 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_27_port, B1 => 
                           n1176, B2 => REGISTERS_21_27_port, ZN => n1268);
   U928 : INV_X1 port map( A => REGISTERS_23_27_port, ZN => n201);
   U929 : INV_X1 port map( A => REGISTERS_22_27_port, ZN => n200);
   U930 : OAI221_X1 port map( B1 => n203, B2 => n1177, C1 => n204, C2 => n1178,
                           A => n1269, ZN => n1262);
   U931 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_27_port, B1 => 
                           n1181, B2 => REGISTERS_17_27_port, ZN => n1269);
   U932 : INV_X1 port map( A => REGISTERS_19_27_port, ZN => n204);
   U933 : INV_X1 port map( A => REGISTERS_18_27_port, ZN => n203);
   U934 : NOR4_X1 port map( A1 => n1270, A2 => n1271, A3 => n1272, A4 => n1273,
                           ZN => n1260);
   U935 : OAI221_X1 port map( B1 => n210, B2 => n1186, C1 => n211, C2 => n1187,
                           A => n1274, ZN => n1273);
   U936 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_27_port, B1 => 
                           n1190, B2 => REGISTERS_13_27_port, ZN => n1274);
   U937 : INV_X1 port map( A => REGISTERS_15_27_port, ZN => n211);
   U938 : INV_X1 port map( A => REGISTERS_14_27_port, ZN => n210);
   U939 : OAI221_X1 port map( B1 => n213, B2 => n1191, C1 => n214, C2 => n1192,
                           A => n1275, ZN => n1272);
   U940 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_27_port, B1 => 
                           n1195, B2 => REGISTERS_9_27_port, ZN => n1275);
   U941 : INV_X1 port map( A => REGISTERS_11_27_port, ZN => n214);
   U942 : INV_X1 port map( A => REGISTERS_10_27_port, ZN => n213);
   U943 : OAI221_X1 port map( B1 => n216, B2 => n1196, C1 => n217, C2 => n1197,
                           A => n1276, ZN => n1271);
   U944 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_27_port, B1 => 
                           n1200, B2 => REGISTERS_5_27_port, ZN => n1276);
   U945 : INV_X1 port map( A => REGISTERS_7_27_port, ZN => n217);
   U946 : INV_X1 port map( A => REGISTERS_6_27_port, ZN => n216);
   U947 : OAI221_X1 port map( B1 => n219, B2 => n1201, C1 => n220, C2 => n1202,
                           A => n1277, ZN => n1270);
   U948 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_27_port, B1 => 
                           n1205, B2 => REGISTERS_1_27_port, ZN => n1277);
   U949 : INV_X1 port map( A => REGISTERS_3_27_port, ZN => n220);
   U950 : INV_X1 port map( A => REGISTERS_2_27_port, ZN => n219);
   U951 : NAND2_X1 port map( A1 => n1278, A2 => n1279, ZN => N2471);
   U952 : NOR4_X1 port map( A1 => n1280, A2 => n1281, A3 => n1282, A4 => n1283,
                           ZN => n1279);
   U953 : OAI221_X1 port map( B1 => n228, B2 => n1162, C1 => n229, C2 => n1163,
                           A => n1284, ZN => n1283);
   U954 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_26_port, B1 => 
                           n1166, B2 => REGISTERS_29_26_port, ZN => n1284);
   U955 : INV_X1 port map( A => REGISTERS_31_26_port, ZN => n229);
   U956 : INV_X1 port map( A => REGISTERS_30_26_port, ZN => n228);
   U957 : OAI221_X1 port map( B1 => n231, B2 => n1167, C1 => n232, C2 => n1168,
                           A => n1285, ZN => n1282);
   U958 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_26_port, B1 => 
                           n1171, B2 => REGISTERS_25_26_port, ZN => n1285);
   U959 : INV_X1 port map( A => REGISTERS_27_26_port, ZN => n232);
   U960 : INV_X1 port map( A => REGISTERS_26_26_port, ZN => n231);
   U961 : OAI221_X1 port map( B1 => n234, B2 => n1172, C1 => n235, C2 => n1173,
                           A => n1286, ZN => n1281);
   U962 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_26_port, B1 => 
                           n1176, B2 => REGISTERS_21_26_port, ZN => n1286);
   U963 : INV_X1 port map( A => REGISTERS_23_26_port, ZN => n235);
   U964 : INV_X1 port map( A => REGISTERS_22_26_port, ZN => n234);
   U965 : OAI221_X1 port map( B1 => n237, B2 => n1177, C1 => n238, C2 => n1178,
                           A => n1287, ZN => n1280);
   U966 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_26_port, B1 => 
                           n1181, B2 => REGISTERS_17_26_port, ZN => n1287);
   U967 : INV_X1 port map( A => REGISTERS_19_26_port, ZN => n238);
   U968 : INV_X1 port map( A => REGISTERS_18_26_port, ZN => n237);
   U969 : NOR4_X1 port map( A1 => n1288, A2 => n1289, A3 => n1290, A4 => n1291,
                           ZN => n1278);
   U970 : OAI221_X1 port map( B1 => n244, B2 => n1186, C1 => n245, C2 => n1187,
                           A => n1292, ZN => n1291);
   U971 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_26_port, B1 => 
                           n1190, B2 => REGISTERS_13_26_port, ZN => n1292);
   U972 : INV_X1 port map( A => REGISTERS_15_26_port, ZN => n245);
   U973 : INV_X1 port map( A => REGISTERS_14_26_port, ZN => n244);
   U974 : OAI221_X1 port map( B1 => n247, B2 => n1191, C1 => n248, C2 => n1192,
                           A => n1293, ZN => n1290);
   U975 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_26_port, B1 => 
                           n1195, B2 => REGISTERS_9_26_port, ZN => n1293);
   U976 : INV_X1 port map( A => REGISTERS_11_26_port, ZN => n248);
   U977 : INV_X1 port map( A => REGISTERS_10_26_port, ZN => n247);
   U978 : OAI221_X1 port map( B1 => n250, B2 => n1196, C1 => n251, C2 => n1197,
                           A => n1294, ZN => n1289);
   U979 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_26_port, B1 => 
                           n1200, B2 => REGISTERS_5_26_port, ZN => n1294);
   U980 : INV_X1 port map( A => REGISTERS_7_26_port, ZN => n251);
   U981 : INV_X1 port map( A => REGISTERS_6_26_port, ZN => n250);
   U982 : OAI221_X1 port map( B1 => n253, B2 => n1201, C1 => n254, C2 => n1202,
                           A => n1295, ZN => n1288);
   U983 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_26_port, B1 => 
                           n1205, B2 => REGISTERS_1_26_port, ZN => n1295);
   U984 : INV_X1 port map( A => REGISTERS_3_26_port, ZN => n254);
   U985 : INV_X1 port map( A => REGISTERS_2_26_port, ZN => n253);
   U986 : NAND2_X1 port map( A1 => n1296, A2 => n1297, ZN => N2469);
   U987 : NOR4_X1 port map( A1 => n1298, A2 => n1299, A3 => n1300, A4 => n1301,
                           ZN => n1297);
   U988 : OAI221_X1 port map( B1 => n262, B2 => n1162, C1 => n263, C2 => n1163,
                           A => n1302, ZN => n1301);
   U989 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_25_port, B1 => 
                           n1166, B2 => REGISTERS_29_25_port, ZN => n1302);
   U990 : INV_X1 port map( A => REGISTERS_31_25_port, ZN => n263);
   U991 : INV_X1 port map( A => REGISTERS_30_25_port, ZN => n262);
   U992 : OAI221_X1 port map( B1 => n265, B2 => n1167, C1 => n266, C2 => n1168,
                           A => n1303, ZN => n1300);
   U993 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_25_port, B1 => 
                           n1171, B2 => REGISTERS_25_25_port, ZN => n1303);
   U994 : INV_X1 port map( A => REGISTERS_27_25_port, ZN => n266);
   U995 : INV_X1 port map( A => REGISTERS_26_25_port, ZN => n265);
   U996 : OAI221_X1 port map( B1 => n268, B2 => n1172, C1 => n269, C2 => n1173,
                           A => n1304, ZN => n1299);
   U997 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_25_port, B1 => 
                           n1176, B2 => REGISTERS_21_25_port, ZN => n1304);
   U998 : INV_X1 port map( A => REGISTERS_23_25_port, ZN => n269);
   U999 : INV_X1 port map( A => REGISTERS_22_25_port, ZN => n268);
   U1000 : OAI221_X1 port map( B1 => n271, B2 => n1177, C1 => n272, C2 => n1178
                           , A => n1305, ZN => n1298);
   U1001 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_25_port, B1 => 
                           n1181, B2 => REGISTERS_17_25_port, ZN => n1305);
   U1002 : INV_X1 port map( A => REGISTERS_19_25_port, ZN => n272);
   U1003 : INV_X1 port map( A => REGISTERS_18_25_port, ZN => n271);
   U1004 : NOR4_X1 port map( A1 => n1306, A2 => n1307, A3 => n1308, A4 => n1309
                           , ZN => n1296);
   U1005 : OAI221_X1 port map( B1 => n278, B2 => n1186, C1 => n279, C2 => n1187
                           , A => n1310, ZN => n1309);
   U1006 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_25_port, B1 => 
                           n1190, B2 => REGISTERS_13_25_port, ZN => n1310);
   U1007 : INV_X1 port map( A => REGISTERS_15_25_port, ZN => n279);
   U1008 : INV_X1 port map( A => REGISTERS_14_25_port, ZN => n278);
   U1009 : OAI221_X1 port map( B1 => n281, B2 => n1191, C1 => n282, C2 => n1192
                           , A => n1311, ZN => n1308);
   U1010 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_25_port, B1 => 
                           n1195, B2 => REGISTERS_9_25_port, ZN => n1311);
   U1011 : INV_X1 port map( A => REGISTERS_11_25_port, ZN => n282);
   U1012 : INV_X1 port map( A => REGISTERS_10_25_port, ZN => n281);
   U1013 : OAI221_X1 port map( B1 => n284, B2 => n1196, C1 => n285, C2 => n1197
                           , A => n1312, ZN => n1307);
   U1014 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_25_port, B1 => 
                           n1200, B2 => REGISTERS_5_25_port, ZN => n1312);
   U1015 : INV_X1 port map( A => REGISTERS_7_25_port, ZN => n285);
   U1016 : INV_X1 port map( A => REGISTERS_6_25_port, ZN => n284);
   U1017 : OAI221_X1 port map( B1 => n287, B2 => n1201, C1 => n288, C2 => n1202
                           , A => n1313, ZN => n1306);
   U1018 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_25_port, B1 => 
                           n1205, B2 => REGISTERS_1_25_port, ZN => n1313);
   U1019 : INV_X1 port map( A => REGISTERS_3_25_port, ZN => n288);
   U1020 : INV_X1 port map( A => REGISTERS_2_25_port, ZN => n287);
   U1021 : NAND2_X1 port map( A1 => n1314, A2 => n1315, ZN => N2467);
   U1022 : NOR4_X1 port map( A1 => n1316, A2 => n1317, A3 => n1318, A4 => n1319
                           , ZN => n1315);
   U1023 : OAI221_X1 port map( B1 => n296, B2 => n1162, C1 => n297, C2 => n1163
                           , A => n1320, ZN => n1319);
   U1024 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_24_port, B1 => 
                           n1166, B2 => REGISTERS_29_24_port, ZN => n1320);
   U1025 : INV_X1 port map( A => REGISTERS_31_24_port, ZN => n297);
   U1026 : INV_X1 port map( A => REGISTERS_30_24_port, ZN => n296);
   U1027 : OAI221_X1 port map( B1 => n299, B2 => n1167, C1 => n300, C2 => n1168
                           , A => n1321, ZN => n1318);
   U1028 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_24_port, B1 => 
                           n1171, B2 => REGISTERS_25_24_port, ZN => n1321);
   U1029 : INV_X1 port map( A => REGISTERS_27_24_port, ZN => n300);
   U1030 : INV_X1 port map( A => REGISTERS_26_24_port, ZN => n299);
   U1031 : OAI221_X1 port map( B1 => n302, B2 => n1172, C1 => n303, C2 => n1173
                           , A => n1322, ZN => n1317);
   U1032 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_24_port, B1 => 
                           n1176, B2 => REGISTERS_21_24_port, ZN => n1322);
   U1033 : INV_X1 port map( A => REGISTERS_23_24_port, ZN => n303);
   U1034 : INV_X1 port map( A => REGISTERS_22_24_port, ZN => n302);
   U1035 : OAI221_X1 port map( B1 => n305, B2 => n1177, C1 => n306, C2 => n1178
                           , A => n1323, ZN => n1316);
   U1036 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_24_port, B1 => 
                           n1181, B2 => REGISTERS_17_24_port, ZN => n1323);
   U1037 : INV_X1 port map( A => REGISTERS_19_24_port, ZN => n306);
   U1038 : INV_X1 port map( A => REGISTERS_18_24_port, ZN => n305);
   U1039 : NOR4_X1 port map( A1 => n1324, A2 => n1325, A3 => n1326, A4 => n1327
                           , ZN => n1314);
   U1040 : OAI221_X1 port map( B1 => n312, B2 => n1186, C1 => n313, C2 => n1187
                           , A => n1328, ZN => n1327);
   U1041 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_24_port, B1 => 
                           n1190, B2 => REGISTERS_13_24_port, ZN => n1328);
   U1042 : INV_X1 port map( A => REGISTERS_15_24_port, ZN => n313);
   U1043 : INV_X1 port map( A => REGISTERS_14_24_port, ZN => n312);
   U1044 : OAI221_X1 port map( B1 => n315, B2 => n1191, C1 => n316, C2 => n1192
                           , A => n1329, ZN => n1326);
   U1045 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_24_port, B1 => 
                           n1195, B2 => REGISTERS_9_24_port, ZN => n1329);
   U1046 : INV_X1 port map( A => REGISTERS_11_24_port, ZN => n316);
   U1047 : INV_X1 port map( A => REGISTERS_10_24_port, ZN => n315);
   U1048 : OAI221_X1 port map( B1 => n318, B2 => n1196, C1 => n319, C2 => n1197
                           , A => n1330, ZN => n1325);
   U1049 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_24_port, B1 => 
                           n1200, B2 => REGISTERS_5_24_port, ZN => n1330);
   U1050 : INV_X1 port map( A => REGISTERS_7_24_port, ZN => n319);
   U1051 : INV_X1 port map( A => REGISTERS_6_24_port, ZN => n318);
   U1052 : OAI221_X1 port map( B1 => n321, B2 => n1201, C1 => n322, C2 => n1202
                           , A => n1331, ZN => n1324);
   U1053 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_24_port, B1 => 
                           n1205, B2 => REGISTERS_1_24_port, ZN => n1331);
   U1054 : INV_X1 port map( A => REGISTERS_3_24_port, ZN => n322);
   U1055 : INV_X1 port map( A => REGISTERS_2_24_port, ZN => n321);
   U1056 : NAND2_X1 port map( A1 => n1332, A2 => n1333, ZN => N2465);
   U1057 : NOR4_X1 port map( A1 => n1334, A2 => n1335, A3 => n1336, A4 => n1337
                           , ZN => n1333);
   U1058 : OAI221_X1 port map( B1 => n330, B2 => n1162, C1 => n331, C2 => n1163
                           , A => n1338, ZN => n1337);
   U1059 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_23_port, B1 => 
                           n1166, B2 => REGISTERS_29_23_port, ZN => n1338);
   U1060 : INV_X1 port map( A => REGISTERS_31_23_port, ZN => n331);
   U1061 : INV_X1 port map( A => REGISTERS_30_23_port, ZN => n330);
   U1062 : OAI221_X1 port map( B1 => n333, B2 => n1167, C1 => n334, C2 => n1168
                           , A => n1339, ZN => n1336);
   U1063 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_23_port, B1 => 
                           n1171, B2 => REGISTERS_25_23_port, ZN => n1339);
   U1064 : INV_X1 port map( A => REGISTERS_27_23_port, ZN => n334);
   U1065 : INV_X1 port map( A => REGISTERS_26_23_port, ZN => n333);
   U1066 : OAI221_X1 port map( B1 => n336, B2 => n1172, C1 => n337, C2 => n1173
                           , A => n1340, ZN => n1335);
   U1067 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_23_port, B1 => 
                           n1176, B2 => REGISTERS_21_23_port, ZN => n1340);
   U1068 : INV_X1 port map( A => REGISTERS_23_23_port, ZN => n337);
   U1069 : INV_X1 port map( A => REGISTERS_22_23_port, ZN => n336);
   U1070 : OAI221_X1 port map( B1 => n339, B2 => n1177, C1 => n340, C2 => n1178
                           , A => n1341, ZN => n1334);
   U1071 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_23_port, B1 => 
                           n1181, B2 => REGISTERS_17_23_port, ZN => n1341);
   U1072 : INV_X1 port map( A => REGISTERS_19_23_port, ZN => n340);
   U1073 : INV_X1 port map( A => REGISTERS_18_23_port, ZN => n339);
   U1074 : NOR4_X1 port map( A1 => n1342, A2 => n1343, A3 => n1344, A4 => n1345
                           , ZN => n1332);
   U1075 : OAI221_X1 port map( B1 => n346, B2 => n1186, C1 => n347, C2 => n1187
                           , A => n1346, ZN => n1345);
   U1076 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_23_port, B1 => 
                           n1190, B2 => REGISTERS_13_23_port, ZN => n1346);
   U1077 : INV_X1 port map( A => REGISTERS_15_23_port, ZN => n347);
   U1078 : INV_X1 port map( A => REGISTERS_14_23_port, ZN => n346);
   U1079 : OAI221_X1 port map( B1 => n349, B2 => n1191, C1 => n350, C2 => n1192
                           , A => n1347, ZN => n1344);
   U1080 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_23_port, B1 => 
                           n1195, B2 => REGISTERS_9_23_port, ZN => n1347);
   U1081 : INV_X1 port map( A => REGISTERS_11_23_port, ZN => n350);
   U1082 : INV_X1 port map( A => REGISTERS_10_23_port, ZN => n349);
   U1083 : OAI221_X1 port map( B1 => n352, B2 => n1196, C1 => n353, C2 => n1197
                           , A => n1348, ZN => n1343);
   U1084 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_23_port, B1 => 
                           n1200, B2 => REGISTERS_5_23_port, ZN => n1348);
   U1085 : INV_X1 port map( A => REGISTERS_7_23_port, ZN => n353);
   U1086 : INV_X1 port map( A => REGISTERS_6_23_port, ZN => n352);
   U1087 : OAI221_X1 port map( B1 => n355, B2 => n1201, C1 => n356, C2 => n1202
                           , A => n1349, ZN => n1342);
   U1088 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_23_port, B1 => 
                           n1205, B2 => REGISTERS_1_23_port, ZN => n1349);
   U1089 : INV_X1 port map( A => REGISTERS_3_23_port, ZN => n356);
   U1090 : INV_X1 port map( A => REGISTERS_2_23_port, ZN => n355);
   U1091 : NAND2_X1 port map( A1 => n1350, A2 => n1351, ZN => N2463);
   U1092 : NOR4_X1 port map( A1 => n1352, A2 => n1353, A3 => n1354, A4 => n1355
                           , ZN => n1351);
   U1093 : OAI221_X1 port map( B1 => n364, B2 => n1162, C1 => n365, C2 => n1163
                           , A => n1356, ZN => n1355);
   U1094 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_22_port, B1 => 
                           n1166, B2 => REGISTERS_29_22_port, ZN => n1356);
   U1095 : INV_X1 port map( A => REGISTERS_31_22_port, ZN => n365);
   U1096 : INV_X1 port map( A => REGISTERS_30_22_port, ZN => n364);
   U1097 : OAI221_X1 port map( B1 => n367, B2 => n1167, C1 => n368, C2 => n1168
                           , A => n1357, ZN => n1354);
   U1098 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_22_port, B1 => 
                           n1171, B2 => REGISTERS_25_22_port, ZN => n1357);
   U1099 : INV_X1 port map( A => REGISTERS_27_22_port, ZN => n368);
   U1100 : INV_X1 port map( A => REGISTERS_26_22_port, ZN => n367);
   U1101 : OAI221_X1 port map( B1 => n370, B2 => n1172, C1 => n371, C2 => n1173
                           , A => n1358, ZN => n1353);
   U1102 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_22_port, B1 => 
                           n1176, B2 => REGISTERS_21_22_port, ZN => n1358);
   U1103 : INV_X1 port map( A => REGISTERS_23_22_port, ZN => n371);
   U1104 : INV_X1 port map( A => REGISTERS_22_22_port, ZN => n370);
   U1105 : OAI221_X1 port map( B1 => n373, B2 => n1177, C1 => n374, C2 => n1178
                           , A => n1359, ZN => n1352);
   U1106 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_22_port, B1 => 
                           n1181, B2 => REGISTERS_17_22_port, ZN => n1359);
   U1107 : INV_X1 port map( A => REGISTERS_19_22_port, ZN => n374);
   U1108 : INV_X1 port map( A => REGISTERS_18_22_port, ZN => n373);
   U1109 : NOR4_X1 port map( A1 => n1360, A2 => n1361, A3 => n1362, A4 => n1363
                           , ZN => n1350);
   U1110 : OAI221_X1 port map( B1 => n380, B2 => n1186, C1 => n381, C2 => n1187
                           , A => n1364, ZN => n1363);
   U1111 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_22_port, B1 => 
                           n1190, B2 => REGISTERS_13_22_port, ZN => n1364);
   U1112 : INV_X1 port map( A => REGISTERS_15_22_port, ZN => n381);
   U1113 : INV_X1 port map( A => REGISTERS_14_22_port, ZN => n380);
   U1114 : OAI221_X1 port map( B1 => n383, B2 => n1191, C1 => n384, C2 => n1192
                           , A => n1365, ZN => n1362);
   U1115 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_22_port, B1 => 
                           n1195, B2 => REGISTERS_9_22_port, ZN => n1365);
   U1116 : INV_X1 port map( A => REGISTERS_11_22_port, ZN => n384);
   U1117 : INV_X1 port map( A => REGISTERS_10_22_port, ZN => n383);
   U1118 : OAI221_X1 port map( B1 => n386, B2 => n1196, C1 => n387, C2 => n1197
                           , A => n1366, ZN => n1361);
   U1119 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_22_port, B1 => 
                           n1200, B2 => REGISTERS_5_22_port, ZN => n1366);
   U1120 : INV_X1 port map( A => REGISTERS_7_22_port, ZN => n387);
   U1121 : INV_X1 port map( A => REGISTERS_6_22_port, ZN => n386);
   U1122 : OAI221_X1 port map( B1 => n389, B2 => n1201, C1 => n390, C2 => n1202
                           , A => n1367, ZN => n1360);
   U1123 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_22_port, B1 => 
                           n1205, B2 => REGISTERS_1_22_port, ZN => n1367);
   U1124 : INV_X1 port map( A => REGISTERS_3_22_port, ZN => n390);
   U1125 : INV_X1 port map( A => REGISTERS_2_22_port, ZN => n389);
   U1126 : NAND2_X1 port map( A1 => n1368, A2 => n1369, ZN => N2461);
   U1127 : NOR4_X1 port map( A1 => n1370, A2 => n1371, A3 => n1372, A4 => n1373
                           , ZN => n1369);
   U1128 : OAI221_X1 port map( B1 => n398, B2 => n1162, C1 => n399, C2 => n1163
                           , A => n1374, ZN => n1373);
   U1129 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_21_port, B1 => 
                           n1166, B2 => REGISTERS_29_21_port, ZN => n1374);
   U1130 : INV_X1 port map( A => REGISTERS_31_21_port, ZN => n399);
   U1131 : INV_X1 port map( A => REGISTERS_30_21_port, ZN => n398);
   U1132 : OAI221_X1 port map( B1 => n401, B2 => n1167, C1 => n402, C2 => n1168
                           , A => n1375, ZN => n1372);
   U1133 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_21_port, B1 => 
                           n1171, B2 => REGISTERS_25_21_port, ZN => n1375);
   U1134 : INV_X1 port map( A => REGISTERS_27_21_port, ZN => n402);
   U1135 : INV_X1 port map( A => REGISTERS_26_21_port, ZN => n401);
   U1136 : OAI221_X1 port map( B1 => n404, B2 => n1172, C1 => n405, C2 => n1173
                           , A => n1376, ZN => n1371);
   U1137 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_21_port, B1 => 
                           n1176, B2 => REGISTERS_21_21_port, ZN => n1376);
   U1138 : INV_X1 port map( A => REGISTERS_23_21_port, ZN => n405);
   U1139 : INV_X1 port map( A => REGISTERS_22_21_port, ZN => n404);
   U1140 : OAI221_X1 port map( B1 => n407, B2 => n1177, C1 => n408, C2 => n1178
                           , A => n1377, ZN => n1370);
   U1141 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_21_port, B1 => 
                           n1181, B2 => REGISTERS_17_21_port, ZN => n1377);
   U1142 : INV_X1 port map( A => REGISTERS_19_21_port, ZN => n408);
   U1143 : INV_X1 port map( A => REGISTERS_18_21_port, ZN => n407);
   U1144 : NOR4_X1 port map( A1 => n1378, A2 => n1379, A3 => n1380, A4 => n1381
                           , ZN => n1368);
   U1145 : OAI221_X1 port map( B1 => n414, B2 => n1186, C1 => n415, C2 => n1187
                           , A => n1382, ZN => n1381);
   U1146 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_21_port, B1 => 
                           n1190, B2 => REGISTERS_13_21_port, ZN => n1382);
   U1147 : INV_X1 port map( A => REGISTERS_15_21_port, ZN => n415);
   U1148 : INV_X1 port map( A => REGISTERS_14_21_port, ZN => n414);
   U1149 : OAI221_X1 port map( B1 => n417, B2 => n1191, C1 => n418, C2 => n1192
                           , A => n1383, ZN => n1380);
   U1150 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_21_port, B1 => 
                           n1195, B2 => REGISTERS_9_21_port, ZN => n1383);
   U1151 : INV_X1 port map( A => REGISTERS_11_21_port, ZN => n418);
   U1152 : INV_X1 port map( A => REGISTERS_10_21_port, ZN => n417);
   U1153 : OAI221_X1 port map( B1 => n420, B2 => n1196, C1 => n421, C2 => n1197
                           , A => n1384, ZN => n1379);
   U1154 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_21_port, B1 => 
                           n1200, B2 => REGISTERS_5_21_port, ZN => n1384);
   U1155 : INV_X1 port map( A => REGISTERS_7_21_port, ZN => n421);
   U1156 : INV_X1 port map( A => REGISTERS_6_21_port, ZN => n420);
   U1157 : OAI221_X1 port map( B1 => n423, B2 => n1201, C1 => n424, C2 => n1202
                           , A => n1385, ZN => n1378);
   U1158 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_21_port, B1 => 
                           n1205, B2 => REGISTERS_1_21_port, ZN => n1385);
   U1159 : INV_X1 port map( A => REGISTERS_3_21_port, ZN => n424);
   U1160 : INV_X1 port map( A => REGISTERS_2_21_port, ZN => n423);
   U1161 : NAND2_X1 port map( A1 => n1386, A2 => n1387, ZN => N2459);
   U1162 : NOR4_X1 port map( A1 => n1388, A2 => n1389, A3 => n1390, A4 => n1391
                           , ZN => n1387);
   U1163 : OAI221_X1 port map( B1 => n432, B2 => n1162, C1 => n433, C2 => n1163
                           , A => n1392, ZN => n1391);
   U1164 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_20_port, B1 => 
                           n1166, B2 => REGISTERS_29_20_port, ZN => n1392);
   U1165 : INV_X1 port map( A => REGISTERS_31_20_port, ZN => n433);
   U1166 : INV_X1 port map( A => REGISTERS_30_20_port, ZN => n432);
   U1167 : OAI221_X1 port map( B1 => n435, B2 => n1167, C1 => n436, C2 => n1168
                           , A => n1393, ZN => n1390);
   U1168 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_20_port, B1 => 
                           n1171, B2 => REGISTERS_25_20_port, ZN => n1393);
   U1169 : INV_X1 port map( A => REGISTERS_27_20_port, ZN => n436);
   U1170 : INV_X1 port map( A => REGISTERS_26_20_port, ZN => n435);
   U1171 : OAI221_X1 port map( B1 => n438, B2 => n1172, C1 => n439, C2 => n1173
                           , A => n1394, ZN => n1389);
   U1172 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_20_port, B1 => 
                           n1176, B2 => REGISTERS_21_20_port, ZN => n1394);
   U1173 : INV_X1 port map( A => REGISTERS_23_20_port, ZN => n439);
   U1174 : INV_X1 port map( A => REGISTERS_22_20_port, ZN => n438);
   U1175 : OAI221_X1 port map( B1 => n441, B2 => n1177, C1 => n442, C2 => n1178
                           , A => n1395, ZN => n1388);
   U1176 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_20_port, B1 => 
                           n1181, B2 => REGISTERS_17_20_port, ZN => n1395);
   U1177 : INV_X1 port map( A => REGISTERS_19_20_port, ZN => n442);
   U1178 : INV_X1 port map( A => REGISTERS_18_20_port, ZN => n441);
   U1179 : NOR4_X1 port map( A1 => n1396, A2 => n1397, A3 => n1398, A4 => n1399
                           , ZN => n1386);
   U1180 : OAI221_X1 port map( B1 => n448, B2 => n1186, C1 => n449, C2 => n1187
                           , A => n1400, ZN => n1399);
   U1181 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_20_port, B1 => 
                           n1190, B2 => REGISTERS_13_20_port, ZN => n1400);
   U1182 : INV_X1 port map( A => REGISTERS_15_20_port, ZN => n449);
   U1183 : INV_X1 port map( A => REGISTERS_14_20_port, ZN => n448);
   U1184 : OAI221_X1 port map( B1 => n451, B2 => n1191, C1 => n452, C2 => n1192
                           , A => n1401, ZN => n1398);
   U1185 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_20_port, B1 => 
                           n1195, B2 => REGISTERS_9_20_port, ZN => n1401);
   U1186 : INV_X1 port map( A => REGISTERS_11_20_port, ZN => n452);
   U1187 : INV_X1 port map( A => REGISTERS_10_20_port, ZN => n451);
   U1188 : OAI221_X1 port map( B1 => n454, B2 => n1196, C1 => n455, C2 => n1197
                           , A => n1402, ZN => n1397);
   U1189 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_20_port, B1 => 
                           n1200, B2 => REGISTERS_5_20_port, ZN => n1402);
   U1190 : INV_X1 port map( A => REGISTERS_7_20_port, ZN => n455);
   U1191 : INV_X1 port map( A => REGISTERS_6_20_port, ZN => n454);
   U1192 : OAI221_X1 port map( B1 => n457, B2 => n1201, C1 => n458, C2 => n1202
                           , A => n1403, ZN => n1396);
   U1193 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_20_port, B1 => 
                           n1205, B2 => REGISTERS_1_20_port, ZN => n1403);
   U1194 : INV_X1 port map( A => REGISTERS_3_20_port, ZN => n458);
   U1195 : INV_X1 port map( A => REGISTERS_2_20_port, ZN => n457);
   U1196 : NAND2_X1 port map( A1 => n1404, A2 => n1405, ZN => N2457);
   U1197 : NOR4_X1 port map( A1 => n1406, A2 => n1407, A3 => n1408, A4 => n1409
                           , ZN => n1405);
   U1198 : OAI221_X1 port map( B1 => n466, B2 => n1162, C1 => n467, C2 => n1163
                           , A => n1410, ZN => n1409);
   U1199 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_19_port, B1 => 
                           n1166, B2 => REGISTERS_29_19_port, ZN => n1410);
   U1200 : INV_X1 port map( A => REGISTERS_31_19_port, ZN => n467);
   U1201 : INV_X1 port map( A => REGISTERS_30_19_port, ZN => n466);
   U1202 : OAI221_X1 port map( B1 => n469, B2 => n1167, C1 => n470, C2 => n1168
                           , A => n1411, ZN => n1408);
   U1203 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_19_port, B1 => 
                           n1171, B2 => REGISTERS_25_19_port, ZN => n1411);
   U1204 : INV_X1 port map( A => REGISTERS_27_19_port, ZN => n470);
   U1205 : INV_X1 port map( A => REGISTERS_26_19_port, ZN => n469);
   U1206 : OAI221_X1 port map( B1 => n472, B2 => n1172, C1 => n473, C2 => n1173
                           , A => n1412, ZN => n1407);
   U1207 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_19_port, B1 => 
                           n1176, B2 => REGISTERS_21_19_port, ZN => n1412);
   U1208 : INV_X1 port map( A => REGISTERS_23_19_port, ZN => n473);
   U1209 : INV_X1 port map( A => REGISTERS_22_19_port, ZN => n472);
   U1210 : OAI221_X1 port map( B1 => n475, B2 => n1177, C1 => n476, C2 => n1178
                           , A => n1413, ZN => n1406);
   U1211 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_19_port, B1 => 
                           n1181, B2 => REGISTERS_17_19_port, ZN => n1413);
   U1212 : INV_X1 port map( A => REGISTERS_19_19_port, ZN => n476);
   U1213 : INV_X1 port map( A => REGISTERS_18_19_port, ZN => n475);
   U1214 : NOR4_X1 port map( A1 => n1414, A2 => n1415, A3 => n1416, A4 => n1417
                           , ZN => n1404);
   U1215 : OAI221_X1 port map( B1 => n482, B2 => n1186, C1 => n483, C2 => n1187
                           , A => n1418, ZN => n1417);
   U1216 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_19_port, B1 => 
                           n1190, B2 => REGISTERS_13_19_port, ZN => n1418);
   U1217 : INV_X1 port map( A => REGISTERS_15_19_port, ZN => n483);
   U1218 : INV_X1 port map( A => REGISTERS_14_19_port, ZN => n482);
   U1219 : OAI221_X1 port map( B1 => n485, B2 => n1191, C1 => n486, C2 => n1192
                           , A => n1419, ZN => n1416);
   U1220 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_19_port, B1 => 
                           n1195, B2 => REGISTERS_9_19_port, ZN => n1419);
   U1221 : INV_X1 port map( A => REGISTERS_11_19_port, ZN => n486);
   U1222 : INV_X1 port map( A => REGISTERS_10_19_port, ZN => n485);
   U1223 : OAI221_X1 port map( B1 => n488, B2 => n1196, C1 => n489, C2 => n1197
                           , A => n1420, ZN => n1415);
   U1224 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_19_port, B1 => 
                           n1200, B2 => REGISTERS_5_19_port, ZN => n1420);
   U1225 : INV_X1 port map( A => REGISTERS_7_19_port, ZN => n489);
   U1226 : INV_X1 port map( A => REGISTERS_6_19_port, ZN => n488);
   U1227 : OAI221_X1 port map( B1 => n491, B2 => n1201, C1 => n492, C2 => n1202
                           , A => n1421, ZN => n1414);
   U1228 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_19_port, B1 => 
                           n1205, B2 => REGISTERS_1_19_port, ZN => n1421);
   U1229 : INV_X1 port map( A => REGISTERS_3_19_port, ZN => n492);
   U1230 : INV_X1 port map( A => REGISTERS_2_19_port, ZN => n491);
   U1231 : NAND2_X1 port map( A1 => n1422, A2 => n1423, ZN => N2455);
   U1232 : NOR4_X1 port map( A1 => n1424, A2 => n1425, A3 => n1426, A4 => n1427
                           , ZN => n1423);
   U1233 : OAI221_X1 port map( B1 => n500, B2 => n1162, C1 => n501, C2 => n1163
                           , A => n1428, ZN => n1427);
   U1234 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_18_port, B1 => 
                           n1166, B2 => REGISTERS_29_18_port, ZN => n1428);
   U1235 : INV_X1 port map( A => REGISTERS_31_18_port, ZN => n501);
   U1236 : INV_X1 port map( A => REGISTERS_30_18_port, ZN => n500);
   U1237 : OAI221_X1 port map( B1 => n503, B2 => n1167, C1 => n504, C2 => n1168
                           , A => n1429, ZN => n1426);
   U1238 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_18_port, B1 => 
                           n1171, B2 => REGISTERS_25_18_port, ZN => n1429);
   U1239 : INV_X1 port map( A => REGISTERS_27_18_port, ZN => n504);
   U1240 : INV_X1 port map( A => REGISTERS_26_18_port, ZN => n503);
   U1241 : OAI221_X1 port map( B1 => n506, B2 => n1172, C1 => n507, C2 => n1173
                           , A => n1430, ZN => n1425);
   U1242 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_18_port, B1 => 
                           n1176, B2 => REGISTERS_21_18_port, ZN => n1430);
   U1243 : INV_X1 port map( A => REGISTERS_23_18_port, ZN => n507);
   U1244 : INV_X1 port map( A => REGISTERS_22_18_port, ZN => n506);
   U1245 : OAI221_X1 port map( B1 => n509, B2 => n1177, C1 => n510, C2 => n1178
                           , A => n1431, ZN => n1424);
   U1246 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_18_port, B1 => 
                           n1181, B2 => REGISTERS_17_18_port, ZN => n1431);
   U1247 : INV_X1 port map( A => REGISTERS_19_18_port, ZN => n510);
   U1248 : INV_X1 port map( A => REGISTERS_18_18_port, ZN => n509);
   U1249 : NOR4_X1 port map( A1 => n1432, A2 => n1433, A3 => n1434, A4 => n1435
                           , ZN => n1422);
   U1250 : OAI221_X1 port map( B1 => n516, B2 => n1186, C1 => n517, C2 => n1187
                           , A => n1436, ZN => n1435);
   U1251 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_18_port, B1 => 
                           n1190, B2 => REGISTERS_13_18_port, ZN => n1436);
   U1252 : INV_X1 port map( A => REGISTERS_15_18_port, ZN => n517);
   U1253 : INV_X1 port map( A => REGISTERS_14_18_port, ZN => n516);
   U1254 : OAI221_X1 port map( B1 => n519, B2 => n1191, C1 => n520, C2 => n1192
                           , A => n1437, ZN => n1434);
   U1255 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_18_port, B1 => 
                           n1195, B2 => REGISTERS_9_18_port, ZN => n1437);
   U1256 : INV_X1 port map( A => REGISTERS_11_18_port, ZN => n520);
   U1257 : INV_X1 port map( A => REGISTERS_10_18_port, ZN => n519);
   U1258 : OAI221_X1 port map( B1 => n522, B2 => n1196, C1 => n523, C2 => n1197
                           , A => n1438, ZN => n1433);
   U1259 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_18_port, B1 => 
                           n1200, B2 => REGISTERS_5_18_port, ZN => n1438);
   U1260 : INV_X1 port map( A => REGISTERS_7_18_port, ZN => n523);
   U1261 : INV_X1 port map( A => REGISTERS_6_18_port, ZN => n522);
   U1262 : OAI221_X1 port map( B1 => n525, B2 => n1201, C1 => n526, C2 => n1202
                           , A => n1439, ZN => n1432);
   U1263 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_18_port, B1 => 
                           n1205, B2 => REGISTERS_1_18_port, ZN => n1439);
   U1264 : INV_X1 port map( A => REGISTERS_3_18_port, ZN => n526);
   U1265 : INV_X1 port map( A => REGISTERS_2_18_port, ZN => n525);
   U1266 : NAND2_X1 port map( A1 => n1440, A2 => n1441, ZN => N2453);
   U1267 : NOR4_X1 port map( A1 => n1442, A2 => n1443, A3 => n1444, A4 => n1445
                           , ZN => n1441);
   U1268 : OAI221_X1 port map( B1 => n534, B2 => n1162, C1 => n535, C2 => n1163
                           , A => n1446, ZN => n1445);
   U1269 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_17_port, B1 => 
                           n1166, B2 => REGISTERS_29_17_port, ZN => n1446);
   U1270 : INV_X1 port map( A => REGISTERS_31_17_port, ZN => n535);
   U1271 : INV_X1 port map( A => REGISTERS_30_17_port, ZN => n534);
   U1272 : OAI221_X1 port map( B1 => n537, B2 => n1167, C1 => n538, C2 => n1168
                           , A => n1447, ZN => n1444);
   U1273 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_17_port, B1 => 
                           n1171, B2 => REGISTERS_25_17_port, ZN => n1447);
   U1274 : INV_X1 port map( A => REGISTERS_27_17_port, ZN => n538);
   U1275 : INV_X1 port map( A => REGISTERS_26_17_port, ZN => n537);
   U1276 : OAI221_X1 port map( B1 => n540, B2 => n1172, C1 => n541, C2 => n1173
                           , A => n1448, ZN => n1443);
   U1277 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_17_port, B1 => 
                           n1176, B2 => REGISTERS_21_17_port, ZN => n1448);
   U1278 : INV_X1 port map( A => REGISTERS_23_17_port, ZN => n541);
   U1279 : INV_X1 port map( A => REGISTERS_22_17_port, ZN => n540);
   U1280 : OAI221_X1 port map( B1 => n543, B2 => n1177, C1 => n544, C2 => n1178
                           , A => n1449, ZN => n1442);
   U1281 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_17_port, B1 => 
                           n1181, B2 => REGISTERS_17_17_port, ZN => n1449);
   U1282 : INV_X1 port map( A => REGISTERS_19_17_port, ZN => n544);
   U1283 : INV_X1 port map( A => REGISTERS_18_17_port, ZN => n543);
   U1284 : NOR4_X1 port map( A1 => n1450, A2 => n1451, A3 => n1452, A4 => n1453
                           , ZN => n1440);
   U1285 : OAI221_X1 port map( B1 => n550, B2 => n1186, C1 => n551, C2 => n1187
                           , A => n1454, ZN => n1453);
   U1286 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_17_port, B1 => 
                           n1190, B2 => REGISTERS_13_17_port, ZN => n1454);
   U1287 : INV_X1 port map( A => REGISTERS_15_17_port, ZN => n551);
   U1288 : INV_X1 port map( A => REGISTERS_14_17_port, ZN => n550);
   U1289 : OAI221_X1 port map( B1 => n553, B2 => n1191, C1 => n554, C2 => n1192
                           , A => n1455, ZN => n1452);
   U1290 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_17_port, B1 => 
                           n1195, B2 => REGISTERS_9_17_port, ZN => n1455);
   U1291 : INV_X1 port map( A => REGISTERS_11_17_port, ZN => n554);
   U1292 : INV_X1 port map( A => REGISTERS_10_17_port, ZN => n553);
   U1293 : OAI221_X1 port map( B1 => n556, B2 => n1196, C1 => n557, C2 => n1197
                           , A => n1456, ZN => n1451);
   U1294 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_17_port, B1 => 
                           n1200, B2 => REGISTERS_5_17_port, ZN => n1456);
   U1295 : INV_X1 port map( A => REGISTERS_7_17_port, ZN => n557);
   U1296 : INV_X1 port map( A => REGISTERS_6_17_port, ZN => n556);
   U1297 : OAI221_X1 port map( B1 => n559, B2 => n1201, C1 => n560, C2 => n1202
                           , A => n1457, ZN => n1450);
   U1298 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_17_port, B1 => 
                           n1205, B2 => REGISTERS_1_17_port, ZN => n1457);
   U1299 : INV_X1 port map( A => REGISTERS_3_17_port, ZN => n560);
   U1300 : INV_X1 port map( A => REGISTERS_2_17_port, ZN => n559);
   U1301 : NAND2_X1 port map( A1 => n1458, A2 => n1459, ZN => N2451);
   U1302 : NOR4_X1 port map( A1 => n1460, A2 => n1461, A3 => n1462, A4 => n1463
                           , ZN => n1459);
   U1303 : OAI221_X1 port map( B1 => n568, B2 => n1162, C1 => n569, C2 => n1163
                           , A => n1464, ZN => n1463);
   U1304 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_16_port, B1 => 
                           n1166, B2 => REGISTERS_29_16_port, ZN => n1464);
   U1305 : INV_X1 port map( A => REGISTERS_31_16_port, ZN => n569);
   U1306 : INV_X1 port map( A => REGISTERS_30_16_port, ZN => n568);
   U1307 : OAI221_X1 port map( B1 => n571, B2 => n1167, C1 => n572, C2 => n1168
                           , A => n1465, ZN => n1462);
   U1308 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_16_port, B1 => 
                           n1171, B2 => REGISTERS_25_16_port, ZN => n1465);
   U1309 : INV_X1 port map( A => REGISTERS_27_16_port, ZN => n572);
   U1310 : INV_X1 port map( A => REGISTERS_26_16_port, ZN => n571);
   U1311 : OAI221_X1 port map( B1 => n574, B2 => n1172, C1 => n575, C2 => n1173
                           , A => n1466, ZN => n1461);
   U1312 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_16_port, B1 => 
                           n1176, B2 => REGISTERS_21_16_port, ZN => n1466);
   U1313 : INV_X1 port map( A => REGISTERS_23_16_port, ZN => n575);
   U1314 : INV_X1 port map( A => REGISTERS_22_16_port, ZN => n574);
   U1315 : OAI221_X1 port map( B1 => n577, B2 => n1177, C1 => n578, C2 => n1178
                           , A => n1467, ZN => n1460);
   U1316 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_16_port, B1 => 
                           n1181, B2 => REGISTERS_17_16_port, ZN => n1467);
   U1317 : INV_X1 port map( A => REGISTERS_19_16_port, ZN => n578);
   U1318 : INV_X1 port map( A => REGISTERS_18_16_port, ZN => n577);
   U1319 : NOR4_X1 port map( A1 => n1468, A2 => n1469, A3 => n1470, A4 => n1471
                           , ZN => n1458);
   U1320 : OAI221_X1 port map( B1 => n584, B2 => n1186, C1 => n585, C2 => n1187
                           , A => n1472, ZN => n1471);
   U1321 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_16_port, B1 => 
                           n1190, B2 => REGISTERS_13_16_port, ZN => n1472);
   U1322 : INV_X1 port map( A => REGISTERS_15_16_port, ZN => n585);
   U1323 : INV_X1 port map( A => REGISTERS_14_16_port, ZN => n584);
   U1324 : OAI221_X1 port map( B1 => n587, B2 => n1191, C1 => n588, C2 => n1192
                           , A => n1473, ZN => n1470);
   U1325 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_16_port, B1 => 
                           n1195, B2 => REGISTERS_9_16_port, ZN => n1473);
   U1326 : INV_X1 port map( A => REGISTERS_11_16_port, ZN => n588);
   U1327 : INV_X1 port map( A => REGISTERS_10_16_port, ZN => n587);
   U1328 : OAI221_X1 port map( B1 => n590, B2 => n1196, C1 => n591, C2 => n1197
                           , A => n1474, ZN => n1469);
   U1329 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_16_port, B1 => 
                           n1200, B2 => REGISTERS_5_16_port, ZN => n1474);
   U1330 : INV_X1 port map( A => REGISTERS_7_16_port, ZN => n591);
   U1331 : INV_X1 port map( A => REGISTERS_6_16_port, ZN => n590);
   U1332 : OAI221_X1 port map( B1 => n593, B2 => n1201, C1 => n594, C2 => n1202
                           , A => n1475, ZN => n1468);
   U1333 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_16_port, B1 => 
                           n1205, B2 => REGISTERS_1_16_port, ZN => n1475);
   U1334 : INV_X1 port map( A => REGISTERS_3_16_port, ZN => n594);
   U1335 : INV_X1 port map( A => REGISTERS_2_16_port, ZN => n593);
   U1336 : NAND2_X1 port map( A1 => n1476, A2 => n1477, ZN => N2449);
   U1337 : NOR4_X1 port map( A1 => n1478, A2 => n1479, A3 => n1480, A4 => n1481
                           , ZN => n1477);
   U1338 : OAI221_X1 port map( B1 => n602, B2 => n1162, C1 => n603, C2 => n1163
                           , A => n1482, ZN => n1481);
   U1339 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_15_port, B1 => 
                           n1166, B2 => REGISTERS_29_15_port, ZN => n1482);
   U1340 : INV_X1 port map( A => REGISTERS_31_15_port, ZN => n603);
   U1341 : INV_X1 port map( A => REGISTERS_30_15_port, ZN => n602);
   U1342 : OAI221_X1 port map( B1 => n605, B2 => n1167, C1 => n606, C2 => n1168
                           , A => n1483, ZN => n1480);
   U1343 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_15_port, B1 => 
                           n1171, B2 => REGISTERS_25_15_port, ZN => n1483);
   U1344 : INV_X1 port map( A => REGISTERS_27_15_port, ZN => n606);
   U1345 : INV_X1 port map( A => REGISTERS_26_15_port, ZN => n605);
   U1346 : OAI221_X1 port map( B1 => n608, B2 => n1172, C1 => n609, C2 => n1173
                           , A => n1484, ZN => n1479);
   U1347 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_15_port, B1 => 
                           n1176, B2 => REGISTERS_21_15_port, ZN => n1484);
   U1348 : INV_X1 port map( A => REGISTERS_23_15_port, ZN => n609);
   U1349 : INV_X1 port map( A => REGISTERS_22_15_port, ZN => n608);
   U1350 : OAI221_X1 port map( B1 => n611, B2 => n1177, C1 => n612, C2 => n1178
                           , A => n1485, ZN => n1478);
   U1351 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_15_port, B1 => 
                           n1181, B2 => REGISTERS_17_15_port, ZN => n1485);
   U1352 : INV_X1 port map( A => REGISTERS_19_15_port, ZN => n612);
   U1353 : INV_X1 port map( A => REGISTERS_18_15_port, ZN => n611);
   U1354 : NOR4_X1 port map( A1 => n1486, A2 => n1487, A3 => n1488, A4 => n1489
                           , ZN => n1476);
   U1355 : OAI221_X1 port map( B1 => n618, B2 => n1186, C1 => n619, C2 => n1187
                           , A => n1490, ZN => n1489);
   U1356 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_15_port, B1 => 
                           n1190, B2 => REGISTERS_13_15_port, ZN => n1490);
   U1357 : INV_X1 port map( A => REGISTERS_15_15_port, ZN => n619);
   U1358 : INV_X1 port map( A => REGISTERS_14_15_port, ZN => n618);
   U1359 : OAI221_X1 port map( B1 => n621, B2 => n1191, C1 => n622, C2 => n1192
                           , A => n1491, ZN => n1488);
   U1360 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_15_port, B1 => 
                           n1195, B2 => REGISTERS_9_15_port, ZN => n1491);
   U1361 : INV_X1 port map( A => REGISTERS_11_15_port, ZN => n622);
   U1362 : INV_X1 port map( A => REGISTERS_10_15_port, ZN => n621);
   U1363 : OAI221_X1 port map( B1 => n624, B2 => n1196, C1 => n625, C2 => n1197
                           , A => n1492, ZN => n1487);
   U1364 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_15_port, B1 => 
                           n1200, B2 => REGISTERS_5_15_port, ZN => n1492);
   U1365 : INV_X1 port map( A => REGISTERS_7_15_port, ZN => n625);
   U1366 : INV_X1 port map( A => REGISTERS_6_15_port, ZN => n624);
   U1367 : OAI221_X1 port map( B1 => n627, B2 => n1201, C1 => n628, C2 => n1202
                           , A => n1493, ZN => n1486);
   U1368 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_15_port, B1 => 
                           n1205, B2 => REGISTERS_1_15_port, ZN => n1493);
   U1369 : INV_X1 port map( A => REGISTERS_3_15_port, ZN => n628);
   U1370 : INV_X1 port map( A => REGISTERS_2_15_port, ZN => n627);
   U1371 : NAND2_X1 port map( A1 => n1494, A2 => n1495, ZN => N2447);
   U1372 : NOR4_X1 port map( A1 => n1496, A2 => n1497, A3 => n1498, A4 => n1499
                           , ZN => n1495);
   U1373 : OAI221_X1 port map( B1 => n636, B2 => n1162, C1 => n637, C2 => n1163
                           , A => n1500, ZN => n1499);
   U1374 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_14_port, B1 => 
                           n1166, B2 => REGISTERS_29_14_port, ZN => n1500);
   U1375 : INV_X1 port map( A => REGISTERS_31_14_port, ZN => n637);
   U1376 : INV_X1 port map( A => REGISTERS_30_14_port, ZN => n636);
   U1377 : OAI221_X1 port map( B1 => n639, B2 => n1167, C1 => n640, C2 => n1168
                           , A => n1501, ZN => n1498);
   U1378 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_14_port, B1 => 
                           n1171, B2 => REGISTERS_25_14_port, ZN => n1501);
   U1379 : INV_X1 port map( A => REGISTERS_27_14_port, ZN => n640);
   U1380 : INV_X1 port map( A => REGISTERS_26_14_port, ZN => n639);
   U1381 : OAI221_X1 port map( B1 => n642, B2 => n1172, C1 => n643, C2 => n1173
                           , A => n1502, ZN => n1497);
   U1382 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_14_port, B1 => 
                           n1176, B2 => REGISTERS_21_14_port, ZN => n1502);
   U1383 : INV_X1 port map( A => REGISTERS_23_14_port, ZN => n643);
   U1384 : INV_X1 port map( A => REGISTERS_22_14_port, ZN => n642);
   U1385 : OAI221_X1 port map( B1 => n645, B2 => n1177, C1 => n646, C2 => n1178
                           , A => n1503, ZN => n1496);
   U1386 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_14_port, B1 => 
                           n1181, B2 => REGISTERS_17_14_port, ZN => n1503);
   U1387 : INV_X1 port map( A => REGISTERS_19_14_port, ZN => n646);
   U1388 : INV_X1 port map( A => REGISTERS_18_14_port, ZN => n645);
   U1389 : NOR4_X1 port map( A1 => n1504, A2 => n1505, A3 => n1506, A4 => n1507
                           , ZN => n1494);
   U1390 : OAI221_X1 port map( B1 => n652, B2 => n1186, C1 => n653, C2 => n1187
                           , A => n1508, ZN => n1507);
   U1391 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_14_port, B1 => 
                           n1190, B2 => REGISTERS_13_14_port, ZN => n1508);
   U1392 : INV_X1 port map( A => REGISTERS_15_14_port, ZN => n653);
   U1393 : INV_X1 port map( A => REGISTERS_14_14_port, ZN => n652);
   U1394 : OAI221_X1 port map( B1 => n655, B2 => n1191, C1 => n656, C2 => n1192
                           , A => n1509, ZN => n1506);
   U1395 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_14_port, B1 => 
                           n1195, B2 => REGISTERS_9_14_port, ZN => n1509);
   U1396 : INV_X1 port map( A => REGISTERS_11_14_port, ZN => n656);
   U1397 : INV_X1 port map( A => REGISTERS_10_14_port, ZN => n655);
   U1398 : OAI221_X1 port map( B1 => n658, B2 => n1196, C1 => n659, C2 => n1197
                           , A => n1510, ZN => n1505);
   U1399 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_14_port, B1 => 
                           n1200, B2 => REGISTERS_5_14_port, ZN => n1510);
   U1400 : INV_X1 port map( A => REGISTERS_7_14_port, ZN => n659);
   U1401 : INV_X1 port map( A => REGISTERS_6_14_port, ZN => n658);
   U1402 : OAI221_X1 port map( B1 => n661, B2 => n1201, C1 => n662, C2 => n1202
                           , A => n1511, ZN => n1504);
   U1403 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_14_port, B1 => 
                           n1205, B2 => REGISTERS_1_14_port, ZN => n1511);
   U1404 : INV_X1 port map( A => REGISTERS_3_14_port, ZN => n662);
   U1405 : INV_X1 port map( A => REGISTERS_2_14_port, ZN => n661);
   U1406 : NAND2_X1 port map( A1 => n1512, A2 => n1513, ZN => N2445);
   U1407 : NOR4_X1 port map( A1 => n1514, A2 => n1515, A3 => n1516, A4 => n1517
                           , ZN => n1513);
   U1408 : OAI221_X1 port map( B1 => n670, B2 => n1162, C1 => n671, C2 => n1163
                           , A => n1518, ZN => n1517);
   U1409 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_13_port, B1 => 
                           n1166, B2 => REGISTERS_29_13_port, ZN => n1518);
   U1410 : INV_X1 port map( A => REGISTERS_31_13_port, ZN => n671);
   U1411 : INV_X1 port map( A => REGISTERS_30_13_port, ZN => n670);
   U1412 : OAI221_X1 port map( B1 => n673, B2 => n1167, C1 => n674, C2 => n1168
                           , A => n1519, ZN => n1516);
   U1413 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_13_port, B1 => 
                           n1171, B2 => REGISTERS_25_13_port, ZN => n1519);
   U1414 : INV_X1 port map( A => REGISTERS_27_13_port, ZN => n674);
   U1415 : INV_X1 port map( A => REGISTERS_26_13_port, ZN => n673);
   U1416 : OAI221_X1 port map( B1 => n676, B2 => n1172, C1 => n677, C2 => n1173
                           , A => n1520, ZN => n1515);
   U1417 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_13_port, B1 => 
                           n1176, B2 => REGISTERS_21_13_port, ZN => n1520);
   U1418 : INV_X1 port map( A => REGISTERS_23_13_port, ZN => n677);
   U1419 : INV_X1 port map( A => REGISTERS_22_13_port, ZN => n676);
   U1420 : OAI221_X1 port map( B1 => n679, B2 => n1177, C1 => n680, C2 => n1178
                           , A => n1521, ZN => n1514);
   U1421 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_13_port, B1 => 
                           n1181, B2 => REGISTERS_17_13_port, ZN => n1521);
   U1422 : INV_X1 port map( A => REGISTERS_19_13_port, ZN => n680);
   U1423 : INV_X1 port map( A => REGISTERS_18_13_port, ZN => n679);
   U1424 : NOR4_X1 port map( A1 => n1522, A2 => n1523, A3 => n1524, A4 => n1525
                           , ZN => n1512);
   U1425 : OAI221_X1 port map( B1 => n686, B2 => n1186, C1 => n687, C2 => n1187
                           , A => n1526, ZN => n1525);
   U1426 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_13_port, B1 => 
                           n1190, B2 => REGISTERS_13_13_port, ZN => n1526);
   U1427 : INV_X1 port map( A => REGISTERS_15_13_port, ZN => n687);
   U1428 : INV_X1 port map( A => REGISTERS_14_13_port, ZN => n686);
   U1429 : OAI221_X1 port map( B1 => n689, B2 => n1191, C1 => n690, C2 => n1192
                           , A => n1527, ZN => n1524);
   U1430 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_13_port, B1 => 
                           n1195, B2 => REGISTERS_9_13_port, ZN => n1527);
   U1431 : INV_X1 port map( A => REGISTERS_11_13_port, ZN => n690);
   U1432 : INV_X1 port map( A => REGISTERS_10_13_port, ZN => n689);
   U1433 : OAI221_X1 port map( B1 => n692, B2 => n1196, C1 => n693, C2 => n1197
                           , A => n1528, ZN => n1523);
   U1434 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_13_port, B1 => 
                           n1200, B2 => REGISTERS_5_13_port, ZN => n1528);
   U1435 : INV_X1 port map( A => REGISTERS_7_13_port, ZN => n693);
   U1436 : INV_X1 port map( A => REGISTERS_6_13_port, ZN => n692);
   U1437 : OAI221_X1 port map( B1 => n695, B2 => n1201, C1 => n696, C2 => n1202
                           , A => n1529, ZN => n1522);
   U1438 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_13_port, B1 => 
                           n1205, B2 => REGISTERS_1_13_port, ZN => n1529);
   U1439 : INV_X1 port map( A => REGISTERS_3_13_port, ZN => n696);
   U1440 : INV_X1 port map( A => REGISTERS_2_13_port, ZN => n695);
   U1441 : NAND2_X1 port map( A1 => n1530, A2 => n1531, ZN => N2443);
   U1442 : NOR4_X1 port map( A1 => n1532, A2 => n1533, A3 => n1534, A4 => n1535
                           , ZN => n1531);
   U1443 : OAI221_X1 port map( B1 => n704, B2 => n1162, C1 => n705, C2 => n1163
                           , A => n1536, ZN => n1535);
   U1444 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_12_port, B1 => 
                           n1166, B2 => REGISTERS_29_12_port, ZN => n1536);
   U1445 : INV_X1 port map( A => REGISTERS_31_12_port, ZN => n705);
   U1446 : INV_X1 port map( A => REGISTERS_30_12_port, ZN => n704);
   U1447 : OAI221_X1 port map( B1 => n707, B2 => n1167, C1 => n708, C2 => n1168
                           , A => n1537, ZN => n1534);
   U1448 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_12_port, B1 => 
                           n1171, B2 => REGISTERS_25_12_port, ZN => n1537);
   U1449 : INV_X1 port map( A => REGISTERS_27_12_port, ZN => n708);
   U1450 : INV_X1 port map( A => REGISTERS_26_12_port, ZN => n707);
   U1451 : OAI221_X1 port map( B1 => n710, B2 => n1172, C1 => n711, C2 => n1173
                           , A => n1538, ZN => n1533);
   U1452 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_12_port, B1 => 
                           n1176, B2 => REGISTERS_21_12_port, ZN => n1538);
   U1453 : INV_X1 port map( A => REGISTERS_23_12_port, ZN => n711);
   U1454 : INV_X1 port map( A => REGISTERS_22_12_port, ZN => n710);
   U1455 : OAI221_X1 port map( B1 => n713, B2 => n1177, C1 => n714, C2 => n1178
                           , A => n1539, ZN => n1532);
   U1456 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_12_port, B1 => 
                           n1181, B2 => REGISTERS_17_12_port, ZN => n1539);
   U1457 : INV_X1 port map( A => REGISTERS_19_12_port, ZN => n714);
   U1458 : INV_X1 port map( A => REGISTERS_18_12_port, ZN => n713);
   U1459 : NOR4_X1 port map( A1 => n1540, A2 => n1541, A3 => n1542, A4 => n1543
                           , ZN => n1530);
   U1460 : OAI221_X1 port map( B1 => n720, B2 => n1186, C1 => n721, C2 => n1187
                           , A => n1544, ZN => n1543);
   U1461 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_12_port, B1 => 
                           n1190, B2 => REGISTERS_13_12_port, ZN => n1544);
   U1462 : INV_X1 port map( A => REGISTERS_15_12_port, ZN => n721);
   U1463 : INV_X1 port map( A => REGISTERS_14_12_port, ZN => n720);
   U1464 : OAI221_X1 port map( B1 => n723, B2 => n1191, C1 => n724, C2 => n1192
                           , A => n1545, ZN => n1542);
   U1465 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_12_port, B1 => 
                           n1195, B2 => REGISTERS_9_12_port, ZN => n1545);
   U1466 : INV_X1 port map( A => REGISTERS_11_12_port, ZN => n724);
   U1467 : INV_X1 port map( A => REGISTERS_10_12_port, ZN => n723);
   U1468 : OAI221_X1 port map( B1 => n726, B2 => n1196, C1 => n727, C2 => n1197
                           , A => n1546, ZN => n1541);
   U1469 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_12_port, B1 => 
                           n1200, B2 => REGISTERS_5_12_port, ZN => n1546);
   U1470 : INV_X1 port map( A => REGISTERS_7_12_port, ZN => n727);
   U1471 : INV_X1 port map( A => REGISTERS_6_12_port, ZN => n726);
   U1472 : OAI221_X1 port map( B1 => n729, B2 => n1201, C1 => n730, C2 => n1202
                           , A => n1547, ZN => n1540);
   U1473 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_12_port, B1 => 
                           n1205, B2 => REGISTERS_1_12_port, ZN => n1547);
   U1474 : INV_X1 port map( A => REGISTERS_3_12_port, ZN => n730);
   U1475 : INV_X1 port map( A => REGISTERS_2_12_port, ZN => n729);
   U1476 : NAND2_X1 port map( A1 => n1548, A2 => n1549, ZN => N2441);
   U1477 : NOR4_X1 port map( A1 => n1550, A2 => n1551, A3 => n1552, A4 => n1553
                           , ZN => n1549);
   U1478 : OAI221_X1 port map( B1 => n738, B2 => n1162, C1 => n739, C2 => n1163
                           , A => n1554, ZN => n1553);
   U1479 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_11_port, B1 => 
                           n1166, B2 => REGISTERS_29_11_port, ZN => n1554);
   U1480 : INV_X1 port map( A => REGISTERS_31_11_port, ZN => n739);
   U1481 : INV_X1 port map( A => REGISTERS_30_11_port, ZN => n738);
   U1482 : OAI221_X1 port map( B1 => n741, B2 => n1167, C1 => n742, C2 => n1168
                           , A => n1555, ZN => n1552);
   U1483 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_11_port, B1 => 
                           n1171, B2 => REGISTERS_25_11_port, ZN => n1555);
   U1484 : INV_X1 port map( A => REGISTERS_27_11_port, ZN => n742);
   U1485 : INV_X1 port map( A => REGISTERS_26_11_port, ZN => n741);
   U1486 : OAI221_X1 port map( B1 => n744, B2 => n1172, C1 => n745, C2 => n1173
                           , A => n1556, ZN => n1551);
   U1487 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_11_port, B1 => 
                           n1176, B2 => REGISTERS_21_11_port, ZN => n1556);
   U1488 : INV_X1 port map( A => REGISTERS_23_11_port, ZN => n745);
   U1489 : INV_X1 port map( A => REGISTERS_22_11_port, ZN => n744);
   U1490 : OAI221_X1 port map( B1 => n747, B2 => n1177, C1 => n748, C2 => n1178
                           , A => n1557, ZN => n1550);
   U1491 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_11_port, B1 => 
                           n1181, B2 => REGISTERS_17_11_port, ZN => n1557);
   U1492 : INV_X1 port map( A => REGISTERS_19_11_port, ZN => n748);
   U1493 : INV_X1 port map( A => REGISTERS_18_11_port, ZN => n747);
   U1494 : NOR4_X1 port map( A1 => n1558, A2 => n1559, A3 => n1560, A4 => n1561
                           , ZN => n1548);
   U1495 : OAI221_X1 port map( B1 => n754, B2 => n1186, C1 => n755, C2 => n1187
                           , A => n1562, ZN => n1561);
   U1496 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_11_port, B1 => 
                           n1190, B2 => REGISTERS_13_11_port, ZN => n1562);
   U1497 : INV_X1 port map( A => REGISTERS_15_11_port, ZN => n755);
   U1498 : INV_X1 port map( A => REGISTERS_14_11_port, ZN => n754);
   U1499 : OAI221_X1 port map( B1 => n757, B2 => n1191, C1 => n758, C2 => n1192
                           , A => n1563, ZN => n1560);
   U1500 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_11_port, B1 => 
                           n1195, B2 => REGISTERS_9_11_port, ZN => n1563);
   U1501 : INV_X1 port map( A => REGISTERS_11_11_port, ZN => n758);
   U1502 : INV_X1 port map( A => REGISTERS_10_11_port, ZN => n757);
   U1503 : OAI221_X1 port map( B1 => n760, B2 => n1196, C1 => n761, C2 => n1197
                           , A => n1564, ZN => n1559);
   U1504 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_11_port, B1 => 
                           n1200, B2 => REGISTERS_5_11_port, ZN => n1564);
   U1505 : INV_X1 port map( A => REGISTERS_7_11_port, ZN => n761);
   U1506 : INV_X1 port map( A => REGISTERS_6_11_port, ZN => n760);
   U1507 : OAI221_X1 port map( B1 => n763, B2 => n1201, C1 => n764, C2 => n1202
                           , A => n1565, ZN => n1558);
   U1508 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_11_port, B1 => 
                           n1205, B2 => REGISTERS_1_11_port, ZN => n1565);
   U1509 : INV_X1 port map( A => REGISTERS_3_11_port, ZN => n764);
   U1510 : INV_X1 port map( A => REGISTERS_2_11_port, ZN => n763);
   U1511 : NAND2_X1 port map( A1 => n1566, A2 => n1567, ZN => N2439);
   U1512 : NOR4_X1 port map( A1 => n1568, A2 => n1569, A3 => n1570, A4 => n1571
                           , ZN => n1567);
   U1513 : OAI221_X1 port map( B1 => n772, B2 => n1162, C1 => n773, C2 => n1163
                           , A => n1572, ZN => n1571);
   U1514 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_10_port, B1 => 
                           n1166, B2 => REGISTERS_29_10_port, ZN => n1572);
   U1515 : INV_X1 port map( A => REGISTERS_31_10_port, ZN => n773);
   U1516 : INV_X1 port map( A => REGISTERS_30_10_port, ZN => n772);
   U1517 : OAI221_X1 port map( B1 => n775, B2 => n1167, C1 => n776, C2 => n1168
                           , A => n1573, ZN => n1570);
   U1518 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_10_port, B1 => 
                           n1171, B2 => REGISTERS_25_10_port, ZN => n1573);
   U1519 : INV_X1 port map( A => REGISTERS_27_10_port, ZN => n776);
   U1520 : INV_X1 port map( A => REGISTERS_26_10_port, ZN => n775);
   U1521 : OAI221_X1 port map( B1 => n778, B2 => n1172, C1 => n779, C2 => n1173
                           , A => n1574, ZN => n1569);
   U1522 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_10_port, B1 => 
                           n1176, B2 => REGISTERS_21_10_port, ZN => n1574);
   U1523 : INV_X1 port map( A => REGISTERS_23_10_port, ZN => n779);
   U1524 : INV_X1 port map( A => REGISTERS_22_10_port, ZN => n778);
   U1525 : OAI221_X1 port map( B1 => n781, B2 => n1177, C1 => n782, C2 => n1178
                           , A => n1575, ZN => n1568);
   U1526 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_10_port, B1 => 
                           n1181, B2 => REGISTERS_17_10_port, ZN => n1575);
   U1527 : INV_X1 port map( A => REGISTERS_19_10_port, ZN => n782);
   U1528 : INV_X1 port map( A => REGISTERS_18_10_port, ZN => n781);
   U1529 : NOR4_X1 port map( A1 => n1576, A2 => n1577, A3 => n1578, A4 => n1579
                           , ZN => n1566);
   U1530 : OAI221_X1 port map( B1 => n788, B2 => n1186, C1 => n789, C2 => n1187
                           , A => n1580, ZN => n1579);
   U1531 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_10_port, B1 => 
                           n1190, B2 => REGISTERS_13_10_port, ZN => n1580);
   U1532 : INV_X1 port map( A => REGISTERS_15_10_port, ZN => n789);
   U1533 : INV_X1 port map( A => REGISTERS_14_10_port, ZN => n788);
   U1534 : OAI221_X1 port map( B1 => n791, B2 => n1191, C1 => n792, C2 => n1192
                           , A => n1581, ZN => n1578);
   U1535 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_10_port, B1 => 
                           n1195, B2 => REGISTERS_9_10_port, ZN => n1581);
   U1536 : INV_X1 port map( A => REGISTERS_11_10_port, ZN => n792);
   U1537 : INV_X1 port map( A => REGISTERS_10_10_port, ZN => n791);
   U1538 : OAI221_X1 port map( B1 => n794, B2 => n1196, C1 => n795, C2 => n1197
                           , A => n1582, ZN => n1577);
   U1539 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_10_port, B1 => 
                           n1200, B2 => REGISTERS_5_10_port, ZN => n1582);
   U1540 : INV_X1 port map( A => REGISTERS_7_10_port, ZN => n795);
   U1541 : INV_X1 port map( A => REGISTERS_6_10_port, ZN => n794);
   U1542 : OAI221_X1 port map( B1 => n797, B2 => n1201, C1 => n798, C2 => n1202
                           , A => n1583, ZN => n1576);
   U1543 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_10_port, B1 => 
                           n1205, B2 => REGISTERS_1_10_port, ZN => n1583);
   U1544 : INV_X1 port map( A => REGISTERS_3_10_port, ZN => n798);
   U1545 : INV_X1 port map( A => REGISTERS_2_10_port, ZN => n797);
   U1546 : NAND2_X1 port map( A1 => n1584, A2 => n1585, ZN => N2437);
   U1547 : NOR4_X1 port map( A1 => n1586, A2 => n1587, A3 => n1588, A4 => n1589
                           , ZN => n1585);
   U1548 : OAI221_X1 port map( B1 => n806, B2 => n1162, C1 => n807, C2 => n1163
                           , A => n1590, ZN => n1589);
   U1549 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_9_port, B1 => 
                           n1166, B2 => REGISTERS_29_9_port, ZN => n1590);
   U1550 : INV_X1 port map( A => REGISTERS_31_9_port, ZN => n807);
   U1551 : INV_X1 port map( A => REGISTERS_30_9_port, ZN => n806);
   U1552 : OAI221_X1 port map( B1 => n809, B2 => n1167, C1 => n810, C2 => n1168
                           , A => n1591, ZN => n1588);
   U1553 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_9_port, B1 => 
                           n1171, B2 => REGISTERS_25_9_port, ZN => n1591);
   U1554 : INV_X1 port map( A => REGISTERS_27_9_port, ZN => n810);
   U1555 : INV_X1 port map( A => REGISTERS_26_9_port, ZN => n809);
   U1556 : OAI221_X1 port map( B1 => n812, B2 => n1172, C1 => n813, C2 => n1173
                           , A => n1592, ZN => n1587);
   U1557 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_9_port, B1 => 
                           n1176, B2 => REGISTERS_21_9_port, ZN => n1592);
   U1558 : INV_X1 port map( A => REGISTERS_23_9_port, ZN => n813);
   U1559 : INV_X1 port map( A => REGISTERS_22_9_port, ZN => n812);
   U1560 : OAI221_X1 port map( B1 => n815, B2 => n1177, C1 => n816, C2 => n1178
                           , A => n1593, ZN => n1586);
   U1561 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_9_port, B1 => 
                           n1181, B2 => REGISTERS_17_9_port, ZN => n1593);
   U1562 : INV_X1 port map( A => REGISTERS_19_9_port, ZN => n816);
   U1563 : INV_X1 port map( A => REGISTERS_18_9_port, ZN => n815);
   U1564 : NOR4_X1 port map( A1 => n1594, A2 => n1595, A3 => n1596, A4 => n1597
                           , ZN => n1584);
   U1565 : OAI221_X1 port map( B1 => n822, B2 => n1186, C1 => n823, C2 => n1187
                           , A => n1598, ZN => n1597);
   U1566 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_9_port, B1 => 
                           n1190, B2 => REGISTERS_13_9_port, ZN => n1598);
   U1567 : INV_X1 port map( A => REGISTERS_15_9_port, ZN => n823);
   U1568 : INV_X1 port map( A => REGISTERS_14_9_port, ZN => n822);
   U1569 : OAI221_X1 port map( B1 => n825, B2 => n1191, C1 => n826, C2 => n1192
                           , A => n1599, ZN => n1596);
   U1570 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_9_port, B1 => 
                           n1195, B2 => REGISTERS_9_9_port, ZN => n1599);
   U1571 : INV_X1 port map( A => REGISTERS_11_9_port, ZN => n826);
   U1572 : INV_X1 port map( A => REGISTERS_10_9_port, ZN => n825);
   U1573 : OAI221_X1 port map( B1 => n828, B2 => n1196, C1 => n829, C2 => n1197
                           , A => n1600, ZN => n1595);
   U1574 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_9_port, B1 => 
                           n1200, B2 => REGISTERS_5_9_port, ZN => n1600);
   U1575 : INV_X1 port map( A => REGISTERS_7_9_port, ZN => n829);
   U1576 : INV_X1 port map( A => REGISTERS_6_9_port, ZN => n828);
   U1577 : OAI221_X1 port map( B1 => n831, B2 => n1201, C1 => n832, C2 => n1202
                           , A => n1601, ZN => n1594);
   U1578 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_9_port, B1 => 
                           n1205, B2 => REGISTERS_1_9_port, ZN => n1601);
   U1579 : INV_X1 port map( A => REGISTERS_3_9_port, ZN => n832);
   U1580 : INV_X1 port map( A => REGISTERS_2_9_port, ZN => n831);
   U1581 : NAND2_X1 port map( A1 => n1602, A2 => n1603, ZN => N2435);
   U1582 : NOR4_X1 port map( A1 => n1604, A2 => n1605, A3 => n1606, A4 => n1607
                           , ZN => n1603);
   U1583 : OAI221_X1 port map( B1 => n840, B2 => n1162, C1 => n841, C2 => n1163
                           , A => n1608, ZN => n1607);
   U1584 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_8_port, B1 => 
                           n1166, B2 => REGISTERS_29_8_port, ZN => n1608);
   U1585 : INV_X1 port map( A => REGISTERS_31_8_port, ZN => n841);
   U1586 : INV_X1 port map( A => REGISTERS_30_8_port, ZN => n840);
   U1587 : OAI221_X1 port map( B1 => n843, B2 => n1167, C1 => n844, C2 => n1168
                           , A => n1609, ZN => n1606);
   U1588 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_8_port, B1 => 
                           n1171, B2 => REGISTERS_25_8_port, ZN => n1609);
   U1589 : INV_X1 port map( A => REGISTERS_27_8_port, ZN => n844);
   U1590 : INV_X1 port map( A => REGISTERS_26_8_port, ZN => n843);
   U1591 : OAI221_X1 port map( B1 => n846, B2 => n1172, C1 => n847, C2 => n1173
                           , A => n1610, ZN => n1605);
   U1592 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_8_port, B1 => 
                           n1176, B2 => REGISTERS_21_8_port, ZN => n1610);
   U1593 : INV_X1 port map( A => REGISTERS_23_8_port, ZN => n847);
   U1594 : INV_X1 port map( A => REGISTERS_22_8_port, ZN => n846);
   U1595 : OAI221_X1 port map( B1 => n849, B2 => n1177, C1 => n850, C2 => n1178
                           , A => n1611, ZN => n1604);
   U1596 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_8_port, B1 => 
                           n1181, B2 => REGISTERS_17_8_port, ZN => n1611);
   U1597 : INV_X1 port map( A => REGISTERS_19_8_port, ZN => n850);
   U1598 : INV_X1 port map( A => REGISTERS_18_8_port, ZN => n849);
   U1599 : NOR4_X1 port map( A1 => n1612, A2 => n1613, A3 => n1614, A4 => n1615
                           , ZN => n1602);
   U1600 : OAI221_X1 port map( B1 => n856, B2 => n1186, C1 => n857, C2 => n1187
                           , A => n1616, ZN => n1615);
   U1601 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_8_port, B1 => 
                           n1190, B2 => REGISTERS_13_8_port, ZN => n1616);
   U1602 : INV_X1 port map( A => REGISTERS_15_8_port, ZN => n857);
   U1603 : INV_X1 port map( A => REGISTERS_14_8_port, ZN => n856);
   U1604 : OAI221_X1 port map( B1 => n859, B2 => n1191, C1 => n860, C2 => n1192
                           , A => n1617, ZN => n1614);
   U1605 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_8_port, B1 => 
                           n1195, B2 => REGISTERS_9_8_port, ZN => n1617);
   U1606 : INV_X1 port map( A => REGISTERS_11_8_port, ZN => n860);
   U1607 : INV_X1 port map( A => REGISTERS_10_8_port, ZN => n859);
   U1608 : OAI221_X1 port map( B1 => n862, B2 => n1196, C1 => n863, C2 => n1197
                           , A => n1618, ZN => n1613);
   U1609 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_8_port, B1 => 
                           n1200, B2 => REGISTERS_5_8_port, ZN => n1618);
   U1610 : INV_X1 port map( A => REGISTERS_7_8_port, ZN => n863);
   U1611 : INV_X1 port map( A => REGISTERS_6_8_port, ZN => n862);
   U1612 : OAI221_X1 port map( B1 => n865, B2 => n1201, C1 => n866, C2 => n1202
                           , A => n1619, ZN => n1612);
   U1613 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_8_port, B1 => 
                           n1205, B2 => REGISTERS_1_8_port, ZN => n1619);
   U1614 : INV_X1 port map( A => REGISTERS_3_8_port, ZN => n866);
   U1615 : INV_X1 port map( A => REGISTERS_2_8_port, ZN => n865);
   U1616 : NAND2_X1 port map( A1 => n1620, A2 => n1621, ZN => N2433);
   U1617 : NOR4_X1 port map( A1 => n1622, A2 => n1623, A3 => n1624, A4 => n1625
                           , ZN => n1621);
   U1618 : OAI221_X1 port map( B1 => n874, B2 => n1162, C1 => n875, C2 => n1163
                           , A => n1626, ZN => n1625);
   U1619 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_7_port, B1 => 
                           n1166, B2 => REGISTERS_29_7_port, ZN => n1626);
   U1620 : INV_X1 port map( A => REGISTERS_31_7_port, ZN => n875);
   U1621 : INV_X1 port map( A => REGISTERS_30_7_port, ZN => n874);
   U1622 : OAI221_X1 port map( B1 => n877, B2 => n1167, C1 => n878, C2 => n1168
                           , A => n1627, ZN => n1624);
   U1623 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_7_port, B1 => 
                           n1171, B2 => REGISTERS_25_7_port, ZN => n1627);
   U1624 : INV_X1 port map( A => REGISTERS_27_7_port, ZN => n878);
   U1625 : INV_X1 port map( A => REGISTERS_26_7_port, ZN => n877);
   U1626 : OAI221_X1 port map( B1 => n880, B2 => n1172, C1 => n881, C2 => n1173
                           , A => n1628, ZN => n1623);
   U1627 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_7_port, B1 => 
                           n1176, B2 => REGISTERS_21_7_port, ZN => n1628);
   U1628 : INV_X1 port map( A => REGISTERS_23_7_port, ZN => n881);
   U1629 : INV_X1 port map( A => REGISTERS_22_7_port, ZN => n880);
   U1630 : OAI221_X1 port map( B1 => n883, B2 => n1177, C1 => n884, C2 => n1178
                           , A => n1629, ZN => n1622);
   U1631 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_7_port, B1 => 
                           n1181, B2 => REGISTERS_17_7_port, ZN => n1629);
   U1632 : INV_X1 port map( A => REGISTERS_19_7_port, ZN => n884);
   U1633 : INV_X1 port map( A => REGISTERS_18_7_port, ZN => n883);
   U1634 : NOR4_X1 port map( A1 => n1630, A2 => n1631, A3 => n1632, A4 => n1633
                           , ZN => n1620);
   U1635 : OAI221_X1 port map( B1 => n890, B2 => n1186, C1 => n891, C2 => n1187
                           , A => n1634, ZN => n1633);
   U1636 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_7_port, B1 => 
                           n1190, B2 => REGISTERS_13_7_port, ZN => n1634);
   U1637 : INV_X1 port map( A => REGISTERS_15_7_port, ZN => n891);
   U1638 : INV_X1 port map( A => REGISTERS_14_7_port, ZN => n890);
   U1639 : OAI221_X1 port map( B1 => n893, B2 => n1191, C1 => n894, C2 => n1192
                           , A => n1635, ZN => n1632);
   U1640 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_7_port, B1 => 
                           n1195, B2 => REGISTERS_9_7_port, ZN => n1635);
   U1641 : INV_X1 port map( A => REGISTERS_11_7_port, ZN => n894);
   U1642 : INV_X1 port map( A => REGISTERS_10_7_port, ZN => n893);
   U1643 : OAI221_X1 port map( B1 => n896, B2 => n1196, C1 => n897, C2 => n1197
                           , A => n1636, ZN => n1631);
   U1644 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_7_port, B1 => 
                           n1200, B2 => REGISTERS_5_7_port, ZN => n1636);
   U1645 : INV_X1 port map( A => REGISTERS_7_7_port, ZN => n897);
   U1646 : INV_X1 port map( A => REGISTERS_6_7_port, ZN => n896);
   U1647 : OAI221_X1 port map( B1 => n899, B2 => n1201, C1 => n900, C2 => n1202
                           , A => n1637, ZN => n1630);
   U1648 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_7_port, B1 => 
                           n1205, B2 => REGISTERS_1_7_port, ZN => n1637);
   U1649 : INV_X1 port map( A => REGISTERS_3_7_port, ZN => n900);
   U1650 : INV_X1 port map( A => REGISTERS_2_7_port, ZN => n899);
   U1651 : NAND2_X1 port map( A1 => n1638, A2 => n1639, ZN => N2431);
   U1652 : NOR4_X1 port map( A1 => n1640, A2 => n1641, A3 => n1642, A4 => n1643
                           , ZN => n1639);
   U1653 : OAI221_X1 port map( B1 => n908, B2 => n1162, C1 => n909, C2 => n1163
                           , A => n1644, ZN => n1643);
   U1654 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_6_port, B1 => 
                           n1166, B2 => REGISTERS_29_6_port, ZN => n1644);
   U1655 : INV_X1 port map( A => REGISTERS_31_6_port, ZN => n909);
   U1656 : INV_X1 port map( A => REGISTERS_30_6_port, ZN => n908);
   U1657 : OAI221_X1 port map( B1 => n911, B2 => n1167, C1 => n912, C2 => n1168
                           , A => n1645, ZN => n1642);
   U1658 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_6_port, B1 => 
                           n1171, B2 => REGISTERS_25_6_port, ZN => n1645);
   U1659 : INV_X1 port map( A => REGISTERS_27_6_port, ZN => n912);
   U1660 : INV_X1 port map( A => REGISTERS_26_6_port, ZN => n911);
   U1661 : OAI221_X1 port map( B1 => n914, B2 => n1172, C1 => n915, C2 => n1173
                           , A => n1646, ZN => n1641);
   U1662 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_6_port, B1 => 
                           n1176, B2 => REGISTERS_21_6_port, ZN => n1646);
   U1663 : INV_X1 port map( A => REGISTERS_23_6_port, ZN => n915);
   U1664 : INV_X1 port map( A => REGISTERS_22_6_port, ZN => n914);
   U1665 : OAI221_X1 port map( B1 => n917, B2 => n1177, C1 => n918, C2 => n1178
                           , A => n1647, ZN => n1640);
   U1666 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_6_port, B1 => 
                           n1181, B2 => REGISTERS_17_6_port, ZN => n1647);
   U1667 : INV_X1 port map( A => REGISTERS_19_6_port, ZN => n918);
   U1668 : INV_X1 port map( A => REGISTERS_18_6_port, ZN => n917);
   U1669 : NOR4_X1 port map( A1 => n1648, A2 => n1649, A3 => n1650, A4 => n1651
                           , ZN => n1638);
   U1670 : OAI221_X1 port map( B1 => n924, B2 => n1186, C1 => n925, C2 => n1187
                           , A => n1652, ZN => n1651);
   U1671 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_6_port, B1 => 
                           n1190, B2 => REGISTERS_13_6_port, ZN => n1652);
   U1672 : INV_X1 port map( A => REGISTERS_15_6_port, ZN => n925);
   U1673 : INV_X1 port map( A => REGISTERS_14_6_port, ZN => n924);
   U1674 : OAI221_X1 port map( B1 => n927, B2 => n1191, C1 => n928, C2 => n1192
                           , A => n1653, ZN => n1650);
   U1675 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_6_port, B1 => 
                           n1195, B2 => REGISTERS_9_6_port, ZN => n1653);
   U1676 : INV_X1 port map( A => REGISTERS_11_6_port, ZN => n928);
   U1677 : INV_X1 port map( A => REGISTERS_10_6_port, ZN => n927);
   U1678 : OAI221_X1 port map( B1 => n930, B2 => n1196, C1 => n931, C2 => n1197
                           , A => n1654, ZN => n1649);
   U1679 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_6_port, B1 => 
                           n1200, B2 => REGISTERS_5_6_port, ZN => n1654);
   U1680 : INV_X1 port map( A => REGISTERS_7_6_port, ZN => n931);
   U1681 : INV_X1 port map( A => REGISTERS_6_6_port, ZN => n930);
   U1682 : OAI221_X1 port map( B1 => n933, B2 => n1201, C1 => n934, C2 => n1202
                           , A => n1655, ZN => n1648);
   U1683 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_6_port, B1 => 
                           n1205, B2 => REGISTERS_1_6_port, ZN => n1655);
   U1684 : INV_X1 port map( A => REGISTERS_3_6_port, ZN => n934);
   U1685 : INV_X1 port map( A => REGISTERS_2_6_port, ZN => n933);
   U1686 : NAND2_X1 port map( A1 => n1656, A2 => n1657, ZN => N2429);
   U1687 : NOR4_X1 port map( A1 => n1658, A2 => n1659, A3 => n1660, A4 => n1661
                           , ZN => n1657);
   U1688 : OAI221_X1 port map( B1 => n942, B2 => n1162, C1 => n943, C2 => n1163
                           , A => n1662, ZN => n1661);
   U1689 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_5_port, B1 => 
                           n1166, B2 => REGISTERS_29_5_port, ZN => n1662);
   U1690 : INV_X1 port map( A => REGISTERS_31_5_port, ZN => n943);
   U1691 : INV_X1 port map( A => REGISTERS_30_5_port, ZN => n942);
   U1692 : OAI221_X1 port map( B1 => n945, B2 => n1167, C1 => n946, C2 => n1168
                           , A => n1663, ZN => n1660);
   U1693 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_5_port, B1 => 
                           n1171, B2 => REGISTERS_25_5_port, ZN => n1663);
   U1694 : INV_X1 port map( A => REGISTERS_27_5_port, ZN => n946);
   U1695 : INV_X1 port map( A => REGISTERS_26_5_port, ZN => n945);
   U1696 : OAI221_X1 port map( B1 => n948, B2 => n1172, C1 => n949, C2 => n1173
                           , A => n1664, ZN => n1659);
   U1697 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_5_port, B1 => 
                           n1176, B2 => REGISTERS_21_5_port, ZN => n1664);
   U1698 : INV_X1 port map( A => REGISTERS_23_5_port, ZN => n949);
   U1699 : INV_X1 port map( A => REGISTERS_22_5_port, ZN => n948);
   U1700 : OAI221_X1 port map( B1 => n951, B2 => n1177, C1 => n952, C2 => n1178
                           , A => n1665, ZN => n1658);
   U1701 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_5_port, B1 => 
                           n1181, B2 => REGISTERS_17_5_port, ZN => n1665);
   U1702 : INV_X1 port map( A => REGISTERS_19_5_port, ZN => n952);
   U1703 : INV_X1 port map( A => REGISTERS_18_5_port, ZN => n951);
   U1704 : NOR4_X1 port map( A1 => n1666, A2 => n1667, A3 => n1668, A4 => n1669
                           , ZN => n1656);
   U1705 : OAI221_X1 port map( B1 => n958, B2 => n1186, C1 => n959, C2 => n1187
                           , A => n1670, ZN => n1669);
   U1706 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_5_port, B1 => 
                           n1190, B2 => REGISTERS_13_5_port, ZN => n1670);
   U1707 : INV_X1 port map( A => REGISTERS_15_5_port, ZN => n959);
   U1708 : INV_X1 port map( A => REGISTERS_14_5_port, ZN => n958);
   U1709 : OAI221_X1 port map( B1 => n961, B2 => n1191, C1 => n962, C2 => n1192
                           , A => n1671, ZN => n1668);
   U1710 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_5_port, B1 => 
                           n1195, B2 => REGISTERS_9_5_port, ZN => n1671);
   U1711 : INV_X1 port map( A => REGISTERS_11_5_port, ZN => n962);
   U1712 : INV_X1 port map( A => REGISTERS_10_5_port, ZN => n961);
   U1713 : OAI221_X1 port map( B1 => n964, B2 => n1196, C1 => n965, C2 => n1197
                           , A => n1672, ZN => n1667);
   U1714 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_5_port, B1 => 
                           n1200, B2 => REGISTERS_5_5_port, ZN => n1672);
   U1715 : INV_X1 port map( A => REGISTERS_7_5_port, ZN => n965);
   U1716 : INV_X1 port map( A => REGISTERS_6_5_port, ZN => n964);
   U1717 : OAI221_X1 port map( B1 => n967, B2 => n1201, C1 => n968, C2 => n1202
                           , A => n1673, ZN => n1666);
   U1718 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_5_port, B1 => 
                           n1205, B2 => REGISTERS_1_5_port, ZN => n1673);
   U1719 : INV_X1 port map( A => REGISTERS_3_5_port, ZN => n968);
   U1720 : INV_X1 port map( A => REGISTERS_2_5_port, ZN => n967);
   U1721 : NAND2_X1 port map( A1 => n1674, A2 => n1675, ZN => N2427);
   U1722 : NOR4_X1 port map( A1 => n1676, A2 => n1677, A3 => n1678, A4 => n1679
                           , ZN => n1675);
   U1723 : OAI221_X1 port map( B1 => n976, B2 => n1162, C1 => n977, C2 => n1163
                           , A => n1680, ZN => n1679);
   U1724 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_4_port, B1 => 
                           n1166, B2 => REGISTERS_29_4_port, ZN => n1680);
   U1725 : INV_X1 port map( A => REGISTERS_31_4_port, ZN => n977);
   U1726 : INV_X1 port map( A => REGISTERS_30_4_port, ZN => n976);
   U1727 : OAI221_X1 port map( B1 => n979, B2 => n1167, C1 => n980, C2 => n1168
                           , A => n1681, ZN => n1678);
   U1728 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_4_port, B1 => 
                           n1171, B2 => REGISTERS_25_4_port, ZN => n1681);
   U1729 : INV_X1 port map( A => REGISTERS_27_4_port, ZN => n980);
   U1730 : INV_X1 port map( A => REGISTERS_26_4_port, ZN => n979);
   U1731 : OAI221_X1 port map( B1 => n982, B2 => n1172, C1 => n983, C2 => n1173
                           , A => n1682, ZN => n1677);
   U1732 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_4_port, B1 => 
                           n1176, B2 => REGISTERS_21_4_port, ZN => n1682);
   U1733 : INV_X1 port map( A => REGISTERS_23_4_port, ZN => n983);
   U1734 : INV_X1 port map( A => REGISTERS_22_4_port, ZN => n982);
   U1735 : OAI221_X1 port map( B1 => n985, B2 => n1177, C1 => n986, C2 => n1178
                           , A => n1683, ZN => n1676);
   U1736 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_4_port, B1 => 
                           n1181, B2 => REGISTERS_17_4_port, ZN => n1683);
   U1737 : INV_X1 port map( A => REGISTERS_19_4_port, ZN => n986);
   U1738 : INV_X1 port map( A => REGISTERS_18_4_port, ZN => n985);
   U1739 : NOR4_X1 port map( A1 => n1684, A2 => n1685, A3 => n1686, A4 => n1687
                           , ZN => n1674);
   U1740 : OAI221_X1 port map( B1 => n992, B2 => n1186, C1 => n993, C2 => n1187
                           , A => n1688, ZN => n1687);
   U1741 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_4_port, B1 => 
                           n1190, B2 => REGISTERS_13_4_port, ZN => n1688);
   U1742 : INV_X1 port map( A => REGISTERS_15_4_port, ZN => n993);
   U1743 : INV_X1 port map( A => REGISTERS_14_4_port, ZN => n992);
   U1744 : OAI221_X1 port map( B1 => n995, B2 => n1191, C1 => n996, C2 => n1192
                           , A => n1689, ZN => n1686);
   U1745 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_4_port, B1 => 
                           n1195, B2 => REGISTERS_9_4_port, ZN => n1689);
   U1746 : INV_X1 port map( A => REGISTERS_11_4_port, ZN => n996);
   U1747 : INV_X1 port map( A => REGISTERS_10_4_port, ZN => n995);
   U1748 : OAI221_X1 port map( B1 => n998, B2 => n1196, C1 => n999, C2 => n1197
                           , A => n1690, ZN => n1685);
   U1749 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_4_port, B1 => 
                           n1200, B2 => REGISTERS_5_4_port, ZN => n1690);
   U1750 : INV_X1 port map( A => REGISTERS_7_4_port, ZN => n999);
   U1751 : INV_X1 port map( A => REGISTERS_6_4_port, ZN => n998);
   U1752 : OAI221_X1 port map( B1 => n1001, B2 => n1201, C1 => n1002, C2 => 
                           n1202, A => n1691, ZN => n1684);
   U1753 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_4_port, B1 => 
                           n1205, B2 => REGISTERS_1_4_port, ZN => n1691);
   U1754 : INV_X1 port map( A => REGISTERS_3_4_port, ZN => n1002);
   U1755 : INV_X1 port map( A => REGISTERS_2_4_port, ZN => n1001);
   U1756 : NAND2_X1 port map( A1 => n1692, A2 => n1693, ZN => N2425);
   U1757 : NOR4_X1 port map( A1 => n1694, A2 => n1695, A3 => n1696, A4 => n1697
                           , ZN => n1693);
   U1758 : OAI221_X1 port map( B1 => n1010, B2 => n1162, C1 => n1011, C2 => 
                           n1163, A => n1698, ZN => n1697);
   U1759 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_3_port, B1 => 
                           n1166, B2 => REGISTERS_29_3_port, ZN => n1698);
   U1760 : INV_X1 port map( A => REGISTERS_31_3_port, ZN => n1011);
   U1761 : INV_X1 port map( A => REGISTERS_30_3_port, ZN => n1010);
   U1762 : OAI221_X1 port map( B1 => n1013, B2 => n1167, C1 => n1014, C2 => 
                           n1168, A => n1699, ZN => n1696);
   U1763 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_3_port, B1 => 
                           n1171, B2 => REGISTERS_25_3_port, ZN => n1699);
   U1764 : INV_X1 port map( A => REGISTERS_27_3_port, ZN => n1014);
   U1765 : INV_X1 port map( A => REGISTERS_26_3_port, ZN => n1013);
   U1766 : OAI221_X1 port map( B1 => n1016, B2 => n1172, C1 => n1017, C2 => 
                           n1173, A => n1700, ZN => n1695);
   U1767 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_3_port, B1 => 
                           n1176, B2 => REGISTERS_21_3_port, ZN => n1700);
   U1768 : INV_X1 port map( A => REGISTERS_23_3_port, ZN => n1017);
   U1769 : INV_X1 port map( A => REGISTERS_22_3_port, ZN => n1016);
   U1770 : OAI221_X1 port map( B1 => n1019, B2 => n1177, C1 => n1020, C2 => 
                           n1178, A => n1701, ZN => n1694);
   U1771 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_3_port, B1 => 
                           n1181, B2 => REGISTERS_17_3_port, ZN => n1701);
   U1772 : INV_X1 port map( A => REGISTERS_19_3_port, ZN => n1020);
   U1773 : INV_X1 port map( A => REGISTERS_18_3_port, ZN => n1019);
   U1774 : NOR4_X1 port map( A1 => n1702, A2 => n1703, A3 => n1704, A4 => n1705
                           , ZN => n1692);
   U1775 : OAI221_X1 port map( B1 => n1026, B2 => n1186, C1 => n1027, C2 => 
                           n1187, A => n1706, ZN => n1705);
   U1776 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_3_port, B1 => 
                           n1190, B2 => REGISTERS_13_3_port, ZN => n1706);
   U1777 : INV_X1 port map( A => REGISTERS_15_3_port, ZN => n1027);
   U1778 : INV_X1 port map( A => REGISTERS_14_3_port, ZN => n1026);
   U1779 : OAI221_X1 port map( B1 => n1029, B2 => n1191, C1 => n1030, C2 => 
                           n1192, A => n1707, ZN => n1704);
   U1780 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_3_port, B1 => 
                           n1195, B2 => REGISTERS_9_3_port, ZN => n1707);
   U1781 : INV_X1 port map( A => REGISTERS_11_3_port, ZN => n1030);
   U1782 : INV_X1 port map( A => REGISTERS_10_3_port, ZN => n1029);
   U1783 : OAI221_X1 port map( B1 => n1032, B2 => n1196, C1 => n1033, C2 => 
                           n1197, A => n1708, ZN => n1703);
   U1784 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_3_port, B1 => 
                           n1200, B2 => REGISTERS_5_3_port, ZN => n1708);
   U1785 : INV_X1 port map( A => REGISTERS_7_3_port, ZN => n1033);
   U1786 : INV_X1 port map( A => REGISTERS_6_3_port, ZN => n1032);
   U1787 : OAI221_X1 port map( B1 => n1035, B2 => n1201, C1 => n1036, C2 => 
                           n1202, A => n1709, ZN => n1702);
   U1788 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_3_port, B1 => 
                           n1205, B2 => REGISTERS_1_3_port, ZN => n1709);
   U1789 : INV_X1 port map( A => REGISTERS_3_3_port, ZN => n1036);
   U1790 : INV_X1 port map( A => REGISTERS_2_3_port, ZN => n1035);
   U1791 : NAND2_X1 port map( A1 => n1710, A2 => n1711, ZN => N2423);
   U1792 : NOR4_X1 port map( A1 => n1712, A2 => n1713, A3 => n1714, A4 => n1715
                           , ZN => n1711);
   U1793 : OAI221_X1 port map( B1 => n1044, B2 => n1162, C1 => n1045, C2 => 
                           n1163, A => n1716, ZN => n1715);
   U1794 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_2_port, B1 => 
                           n1166, B2 => REGISTERS_29_2_port, ZN => n1716);
   U1795 : INV_X1 port map( A => REGISTERS_31_2_port, ZN => n1045);
   U1796 : INV_X1 port map( A => REGISTERS_30_2_port, ZN => n1044);
   U1797 : OAI221_X1 port map( B1 => n1047, B2 => n1167, C1 => n1048, C2 => 
                           n1168, A => n1717, ZN => n1714);
   U1798 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_2_port, B1 => 
                           n1171, B2 => REGISTERS_25_2_port, ZN => n1717);
   U1799 : INV_X1 port map( A => REGISTERS_27_2_port, ZN => n1048);
   U1800 : INV_X1 port map( A => REGISTERS_26_2_port, ZN => n1047);
   U1801 : OAI221_X1 port map( B1 => n1050, B2 => n1172, C1 => n1051, C2 => 
                           n1173, A => n1718, ZN => n1713);
   U1802 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_2_port, B1 => 
                           n1176, B2 => REGISTERS_21_2_port, ZN => n1718);
   U1803 : INV_X1 port map( A => REGISTERS_23_2_port, ZN => n1051);
   U1804 : INV_X1 port map( A => REGISTERS_22_2_port, ZN => n1050);
   U1805 : OAI221_X1 port map( B1 => n1053, B2 => n1177, C1 => n1054, C2 => 
                           n1178, A => n1719, ZN => n1712);
   U1806 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_2_port, B1 => 
                           n1181, B2 => REGISTERS_17_2_port, ZN => n1719);
   U1807 : INV_X1 port map( A => REGISTERS_19_2_port, ZN => n1054);
   U1808 : INV_X1 port map( A => REGISTERS_18_2_port, ZN => n1053);
   U1809 : NOR4_X1 port map( A1 => n1720, A2 => n1721, A3 => n1722, A4 => n1723
                           , ZN => n1710);
   U1810 : OAI221_X1 port map( B1 => n1060, B2 => n1186, C1 => n1061, C2 => 
                           n1187, A => n1724, ZN => n1723);
   U1811 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_2_port, B1 => 
                           n1190, B2 => REGISTERS_13_2_port, ZN => n1724);
   U1812 : INV_X1 port map( A => REGISTERS_15_2_port, ZN => n1061);
   U1813 : INV_X1 port map( A => REGISTERS_14_2_port, ZN => n1060);
   U1814 : OAI221_X1 port map( B1 => n1063, B2 => n1191, C1 => n1064, C2 => 
                           n1192, A => n1725, ZN => n1722);
   U1815 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_2_port, B1 => 
                           n1195, B2 => REGISTERS_9_2_port, ZN => n1725);
   U1816 : INV_X1 port map( A => REGISTERS_11_2_port, ZN => n1064);
   U1817 : INV_X1 port map( A => REGISTERS_10_2_port, ZN => n1063);
   U1818 : OAI221_X1 port map( B1 => n1066, B2 => n1196, C1 => n1067, C2 => 
                           n1197, A => n1726, ZN => n1721);
   U1819 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_2_port, B1 => 
                           n1200, B2 => REGISTERS_5_2_port, ZN => n1726);
   U1820 : INV_X1 port map( A => REGISTERS_7_2_port, ZN => n1067);
   U1821 : INV_X1 port map( A => REGISTERS_6_2_port, ZN => n1066);
   U1822 : OAI221_X1 port map( B1 => n1069, B2 => n1201, C1 => n1070, C2 => 
                           n1202, A => n1727, ZN => n1720);
   U1823 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_2_port, B1 => 
                           n1205, B2 => REGISTERS_1_2_port, ZN => n1727);
   U1824 : INV_X1 port map( A => REGISTERS_3_2_port, ZN => n1070);
   U1825 : INV_X1 port map( A => REGISTERS_2_2_port, ZN => n1069);
   U1826 : NAND2_X1 port map( A1 => n1728, A2 => n1729, ZN => N2421);
   U1827 : NOR4_X1 port map( A1 => n1730, A2 => n1731, A3 => n1732, A4 => n1733
                           , ZN => n1729);
   U1828 : OAI221_X1 port map( B1 => n1078, B2 => n1162, C1 => n1079, C2 => 
                           n1163, A => n1734, ZN => n1733);
   U1829 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_1_port, B1 => 
                           n1166, B2 => REGISTERS_29_1_port, ZN => n1734);
   U1830 : INV_X1 port map( A => REGISTERS_31_1_port, ZN => n1079);
   U1831 : INV_X1 port map( A => REGISTERS_30_1_port, ZN => n1078);
   U1832 : OAI221_X1 port map( B1 => n1081, B2 => n1167, C1 => n1082, C2 => 
                           n1168, A => n1735, ZN => n1732);
   U1833 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_1_port, B1 => 
                           n1171, B2 => REGISTERS_25_1_port, ZN => n1735);
   U1834 : INV_X1 port map( A => REGISTERS_27_1_port, ZN => n1082);
   U1835 : INV_X1 port map( A => REGISTERS_26_1_port, ZN => n1081);
   U1836 : OAI221_X1 port map( B1 => n1084, B2 => n1172, C1 => n1085, C2 => 
                           n1173, A => n1736, ZN => n1731);
   U1837 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_1_port, B1 => 
                           n1176, B2 => REGISTERS_21_1_port, ZN => n1736);
   U1838 : INV_X1 port map( A => REGISTERS_23_1_port, ZN => n1085);
   U1839 : INV_X1 port map( A => REGISTERS_22_1_port, ZN => n1084);
   U1840 : OAI221_X1 port map( B1 => n1087, B2 => n1177, C1 => n1088, C2 => 
                           n1178, A => n1737, ZN => n1730);
   U1841 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_1_port, B1 => 
                           n1181, B2 => REGISTERS_17_1_port, ZN => n1737);
   U1842 : INV_X1 port map( A => REGISTERS_19_1_port, ZN => n1088);
   U1843 : INV_X1 port map( A => REGISTERS_18_1_port, ZN => n1087);
   U1844 : NOR4_X1 port map( A1 => n1738, A2 => n1739, A3 => n1740, A4 => n1741
                           , ZN => n1728);
   U1845 : OAI221_X1 port map( B1 => n1094, B2 => n1186, C1 => n1095, C2 => 
                           n1187, A => n1742, ZN => n1741);
   U1846 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_1_port, B1 => 
                           n1190, B2 => REGISTERS_13_1_port, ZN => n1742);
   U1847 : INV_X1 port map( A => REGISTERS_15_1_port, ZN => n1095);
   U1848 : INV_X1 port map( A => REGISTERS_14_1_port, ZN => n1094);
   U1849 : OAI221_X1 port map( B1 => n1097, B2 => n1191, C1 => n1098, C2 => 
                           n1192, A => n1743, ZN => n1740);
   U1850 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_1_port, B1 => 
                           n1195, B2 => REGISTERS_9_1_port, ZN => n1743);
   U1851 : INV_X1 port map( A => REGISTERS_11_1_port, ZN => n1098);
   U1852 : INV_X1 port map( A => REGISTERS_10_1_port, ZN => n1097);
   U1853 : OAI221_X1 port map( B1 => n1100, B2 => n1196, C1 => n1101, C2 => 
                           n1197, A => n1744, ZN => n1739);
   U1854 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_1_port, B1 => 
                           n1200, B2 => REGISTERS_5_1_port, ZN => n1744);
   U1855 : INV_X1 port map( A => REGISTERS_7_1_port, ZN => n1101);
   U1856 : INV_X1 port map( A => REGISTERS_6_1_port, ZN => n1100);
   U1857 : OAI221_X1 port map( B1 => n1103, B2 => n1201, C1 => n1104, C2 => 
                           n1202, A => n1745, ZN => n1738);
   U1858 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_1_port, B1 => 
                           n1205, B2 => REGISTERS_1_1_port, ZN => n1745);
   U1859 : INV_X1 port map( A => REGISTERS_3_1_port, ZN => n1104);
   U1860 : INV_X1 port map( A => REGISTERS_2_1_port, ZN => n1103);
   U1861 : NAND2_X1 port map( A1 => n1746, A2 => n1747, ZN => N2419);
   U1862 : NOR4_X1 port map( A1 => n1748, A2 => n1749, A3 => n1750, A4 => n1751
                           , ZN => n1747);
   U1863 : OAI221_X1 port map( B1 => n1112, B2 => n1162, C1 => n1113, C2 => 
                           n1163, A => n1752, ZN => n1751);
   U1864 : AOI22_X1 port map( A1 => n1165, A2 => REGISTERS_28_0_port, B1 => 
                           n1166, B2 => REGISTERS_29_0_port, ZN => n1752);
   U1865 : INV_X1 port map( A => REGISTERS_31_0_port, ZN => n1113);
   U1866 : INV_X1 port map( A => REGISTERS_30_0_port, ZN => n1112);
   U1867 : OAI221_X1 port map( B1 => n1119, B2 => n1167, C1 => n1120, C2 => 
                           n1168, A => n1757, ZN => n1750);
   U1868 : AOI22_X1 port map( A1 => n1170, A2 => REGISTERS_24_0_port, B1 => 
                           n1171, B2 => REGISTERS_25_0_port, ZN => n1757);
   U1869 : AND3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(3), ZN => n1753);
   U1870 : INV_X1 port map( A => REGISTERS_27_0_port, ZN => n1120);
   U1871 : AND3_X1 port map( A1 => ADD_RD1(4), A2 => n1760, A3 => ADD_RD1(3), 
                           ZN => n1755);
   U1872 : INV_X1 port map( A => REGISTERS_26_0_port, ZN => n1119);
   U1873 : OAI221_X1 port map( B1 => n1125, B2 => n1172, C1 => n1126, C2 => 
                           n1173, A => n1761, ZN => n1749);
   U1874 : AOI22_X1 port map( A1 => n1175, A2 => REGISTERS_20_0_port, B1 => 
                           n1176, B2 => REGISTERS_21_0_port, ZN => n1761);
   U1875 : INV_X1 port map( A => REGISTERS_23_0_port, ZN => n1126);
   U1876 : INV_X1 port map( A => REGISTERS_22_0_port, ZN => n1125);
   U1877 : OAI221_X1 port map( B1 => n1130, B2 => n1177, C1 => n1131, C2 => 
                           n1178, A => n1764, ZN => n1748);
   U1878 : AOI22_X1 port map( A1 => n1180, A2 => REGISTERS_16_0_port, B1 => 
                           n1181, B2 => REGISTERS_17_0_port, ZN => n1764);
   U1879 : AND3_X1 port map( A1 => ADD_RD1(4), A2 => n1765, A3 => ADD_RD1(0), 
                           ZN => n1762);
   U1880 : INV_X1 port map( A => REGISTERS_19_0_port, ZN => n1131);
   U1881 : AND3_X1 port map( A1 => n1760, A2 => n1765, A3 => ADD_RD1(4), ZN => 
                           n1763);
   U1882 : INV_X1 port map( A => REGISTERS_18_0_port, ZN => n1130);
   U1883 : NOR4_X1 port map( A1 => n1766, A2 => n1767, A3 => n1768, A4 => n1769
                           , ZN => n1746);
   U1884 : OAI221_X1 port map( B1 => n1138, B2 => n1186, C1 => n1139, C2 => 
                           n1187, A => n1770, ZN => n1769);
   U1885 : AOI22_X1 port map( A1 => n1189, A2 => REGISTERS_12_0_port, B1 => 
                           n1190, B2 => REGISTERS_13_0_port, ZN => n1770);
   U1886 : INV_X1 port map( A => REGISTERS_15_0_port, ZN => n1139);
   U1887 : INV_X1 port map( A => REGISTERS_14_0_port, ZN => n1138);
   U1888 : OAI221_X1 port map( B1 => n1143, B2 => n1191, C1 => n1144, C2 => 
                           n1192, A => n1773, ZN => n1768);
   U1889 : AOI22_X1 port map( A1 => n1194, A2 => REGISTERS_8_0_port, B1 => 
                           n1195, B2 => REGISTERS_9_0_port, ZN => n1773);
   U1890 : NOR3_X1 port map( A1 => n1760, A2 => ADD_RD1(4), A3 => n1765, ZN => 
                           n1771);
   U1891 : INV_X1 port map( A => REGISTERS_11_0_port, ZN => n1144);
   U1892 : NOR3_X1 port map( A1 => ADD_RD1(0), A2 => ADD_RD1(4), A3 => n1765, 
                           ZN => n1772);
   U1893 : INV_X1 port map( A => ADD_RD1(3), ZN => n1765);
   U1894 : INV_X1 port map( A => REGISTERS_10_0_port, ZN => n1143);
   U1895 : OAI221_X1 port map( B1 => n1146, B2 => n1196, C1 => n1147, C2 => 
                           n1197, A => n1774, ZN => n1767);
   U1896 : AOI22_X1 port map( A1 => n1199, A2 => REGISTERS_4_0_port, B1 => 
                           n1200, B2 => REGISTERS_5_0_port, ZN => n1774);
   U1897 : AND3_X1 port map( A1 => n1151, A2 => n1777, A3 => ADD_RD1(2), ZN => 
                           n1754);
   U1898 : INV_X1 port map( A => REGISTERS_7_0_port, ZN => n1147);
   U1899 : AND3_X1 port map( A1 => ADD_RD1(1), A2 => n1151, A3 => ADD_RD1(2), 
                           ZN => n1756);
   U1900 : INV_X1 port map( A => n85, ZN => n1151);
   U1901 : INV_X1 port map( A => REGISTERS_6_0_port, ZN => n1146);
   U1902 : OAI221_X1 port map( B1 => n1153, B2 => n1201, C1 => n1154, C2 => 
                           n1202, A => n1778, ZN => n1766);
   U1903 : AOI22_X1 port map( A1 => n1204, A2 => REGISTERS_0_0_port, B1 => 
                           n1205, B2 => REGISTERS_1_0_port, ZN => n1778);
   U1904 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => n1760, 
                           ZN => n1775);
   U1905 : INV_X1 port map( A => ADD_RD1(0), ZN => n1760);
   U1906 : INV_X1 port map( A => REGISTERS_3_0_port, ZN => n1154);
   U1907 : INV_X1 port map( A => ADD_RD1(1), ZN => n1777);
   U1908 : NAND2_X1 port map( A1 => ENABLE, A2 => RESET, ZN => n85);
   U1909 : NOR3_X1 port map( A1 => ADD_RD1(3), A2 => ADD_RD1(4), A3 => 
                           ADD_RD1(0), ZN => n1776);
   U1910 : INV_X1 port map( A => REGISTERS_2_0_port, ZN => n1153);

end SYN_A;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity 
   CU_HDW_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE21 is

   port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0);  
         flush : in std_logic;  IR_LATCH_EN, NPC1_LATCH_EN, NPC2_LATCH_EN, 
         RegA_LATCH_EN, RegB_LATCH_EN, RegAluOpCodeGen_EN, RegIMM_LATCH_EN, 
         Reg_RD1_EN, RD1, RD2, B2_LATCH_EN, MUXA_SEL, MUXB_SEL, ALU_OUTREG_EN, 
         RETURN_REG_EN, Reg_RD2_EN, DRAM_WE, ALU_OUT2_SEL, LMD_LATCH_EN, 
         Alu_outreg2_en, JUMP_en, PC_LATCH_EN, Reg_RD3_EN, write_stop_if_branch
         , WB_MUX_SEL, RF_WE, WB_MUX_ADD_SEL, WR : out std_logic);

end CU_HDW_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE21;

architecture SYN_beh of 
   CU_HDW_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NOR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI211_X1
      port( C1, C2, A, B : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OAI21_X1
      port( B1, B2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component OR4_X1
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component AOI221_X1
      port( B1, B2, C1, C2, A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X8
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X4
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFR_X2
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFF_X1
      port( D, CK : in std_logic;  Q, QN : out std_logic);
   end component;
   
   component DFFS_X1
      port( D, CK, SN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal IR_LATCH_EN_port, RD1_port, RD2_port, RegAluOpCodeGen_EN_port, 
      RegIMM_LATCH_EN_port, Reg_RD1_EN_port, cw_19_port, cw_18_port, cw_17_port
      , cw_15_port, cw_14_port, cw_9_port, cw_8_port, cw_7_port, cw_6_port, 
      cw_5_port, cw_4_port, cw_2_port, cw1_19_port, cw1_18_port, cw1_17_port, 
      cw1_16_port, cw1_15_port, cw1_14_port, cw1_13_port, cw1_12_port, 
      cw1_11_port, cw1_10_port, cw1_9_port, cw1_8_port, cw1_7_port, cw1_6_port,
      cw1_5_port, cw1_4_port, cw1_3_port, cw1_2_port, cw1_1_port, cw1_0_port, 
      cw2_15_port, cw2_14_port, cw2_13_port, cw2_12_port, cw2_11_port, 
      cw2_10_port, cw2_9_port, cw2_8_port, cw2_7_port, cw2_6_port, cw2_5_port, 
      cw2_4_port, cw2_3_port, cw2_2_port, cw2_1_port, cw2_0_port, cw3_10_port, 
      cw3_9_port, cw3_8_port, cw3_7_port, cw3_6_port, cw3_5_port, cw3_4_port, 
      cw3_3_port, cw3_2_port, cw3_1_port, cw3_0_port, cw4_3_port, cw4_2_port, 
      cw4_1_port, cw4_0_port, N442, n37, n38, n39, n42, n43, n44, n45, n48, n49
      , n50, n51, n54, n56, n57, n60, n61, n62, n65, n66, n67, n70, n71, n72, 
      n75, n77, n80, n82, n85, n87, n90, n91, n92, n95, n96, n99, n100, n103, 
      n107, n111, n115, n118, n121, n124, n127, n129, n131, n133, n135, n137, 
      n139, n141, n143, n145, n147, n149, n151, n153, n155, n157, n159, n161, 
      n163, n165, n167, n169, n1, n2, n3, n4, n5, n6, n7, B2_LATCH_EN_port, n9,
      NPC1_LATCH_EN_port, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21
      , n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, 
      n36, n40, n41, n46, n47, n52, n53, n55, n58, net43115, net43116, net43117
      , net43118, net43119, net43120, net43121, net43122, net43123, net43124, 
      net43125, net43126, net43127, net43128, net43129, net43130, net43131, 
      net43132, net43133, net43134, net43135, net43136, net43137, net43138, 
      net43139, net43140, net43141, net43142, net43143, net43144, net43145, 
      net43146, net43147, net43148, net43149, net43150, net43151, net43152, 
      net43153, net43154, net43155, net43156, net43157, net43158, net43159, 
      net43160, net43161, net43162, net43163, net43164, net43165, net43166, 
      net43167, net43168, net43169, net43170, net43171, net43172, net43173, 
      net43174, net43175, net43176, net43177, net43178, net43179, net43180, 
      net43181, net43182, net43183, net43184, net43185, net43186, net43187, 
      net43188, net43189, net43190, net43191, net43192, net43193, net43194, 
      net43195, net43196 : std_logic;

begin
   IR_LATCH_EN <= NPC1_LATCH_EN_port;
   NPC1_LATCH_EN <= NPC1_LATCH_EN_port;
   NPC2_LATCH_EN <= RegAluOpCodeGen_EN_port;
   RegA_LATCH_EN <= RD1_port;
   RegB_LATCH_EN <= RD2_port;
   RegAluOpCodeGen_EN <= RegAluOpCodeGen_EN_port;
   RegIMM_LATCH_EN <= RegIMM_LATCH_EN_port;
   Reg_RD1_EN <= Reg_RD1_EN_port;
   RD1 <= RD1_port;
   RD2 <= RD2_port;
   B2_LATCH_EN <= B2_LATCH_EN_port;
   RETURN_REG_EN <= B2_LATCH_EN_port;
   
   cw1_reg_20_inst : DFFS_X1 port map( D => cw_6_port, CK => N442, SN => Rst, Q
                           => IR_LATCH_EN_port, QN => net43196);
   cw1_reg_19_inst : DFFR_X1 port map( D => cw_19_port, CK => N442, RN => Rst, 
                           Q => cw1_19_port, QN => net43195);
   cw1_reg_18_inst : DFFR_X1 port map( D => cw_18_port, CK => N442, RN => Rst, 
                           Q => cw1_18_port, QN => net43194);
   cw1_reg_17_inst : DFFR_X1 port map( D => cw_17_port, CK => N442, RN => Rst, 
                           Q => cw1_17_port, QN => net43193);
   cw1_reg_16_inst : DFFR_X1 port map( D => cw_5_port, CK => N442, RN => Rst, Q
                           => cw1_16_port, QN => net43192);
   cw1_reg_15_inst : DFFR_X1 port map( D => cw_15_port, CK => N442, RN => Rst, 
                           Q => cw1_15_port, QN => net43191);
   cw1_reg_14_inst : DFFR_X1 port map( D => cw_14_port, CK => N442, RN => Rst, 
                           Q => cw1_14_port, QN => net43190);
   cw1_reg_13_inst : DFFR_X1 port map( D => cw_7_port, CK => N442, RN => Rst, Q
                           => cw1_13_port, QN => net43189);
   cw1_reg_12_inst : DFFR_X1 port map( D => cw_5_port, CK => N442, RN => Rst, Q
                           => cw1_12_port, QN => net43188);
   cw1_reg_11_inst : DFFR_X1 port map( D => cw_15_port, CK => N442, RN => Rst, 
                           Q => cw1_11_port, QN => net43187);
   cw1_reg_10_inst : DFFR_X1 port map( D => cw_8_port, CK => N442, RN => Rst, Q
                           => cw1_10_port, QN => net43186);
   cw1_reg_9_inst : DFFR_X1 port map( D => cw_9_port, CK => N442, RN => Rst, Q 
                           => cw1_9_port, QN => net43185);
   cw1_reg_8_inst : DFFR_X1 port map( D => cw_8_port, CK => N442, RN => Rst, Q 
                           => cw1_8_port, QN => net43184);
   cw1_reg_7_inst : DFFR_X1 port map( D => cw_7_port, CK => N442, RN => Rst, Q 
                           => cw1_7_port, QN => net43183);
   cw1_reg_6_inst : DFFR_X1 port map( D => cw_6_port, CK => N442, RN => Rst, Q 
                           => cw1_6_port, QN => net43182);
   cw1_reg_5_inst : DFFR_X1 port map( D => cw_5_port, CK => N442, RN => Rst, Q 
                           => cw1_5_port, QN => net43181);
   cw1_reg_4_inst : DFFR_X1 port map( D => cw_4_port, CK => N442, RN => Rst, Q 
                           => cw1_4_port, QN => net43180);
   cw1_reg_3_inst : DFFR_X1 port map( D => cw_8_port, CK => N442, RN => Rst, Q 
                           => cw1_3_port, QN => net43179);
   cw1_reg_2_inst : DFFR_X1 port map( D => cw_2_port, CK => N442, RN => Rst, Q 
                           => cw1_2_port, QN => net43178);
   cw1_reg_1_inst : DFFR_X1 port map( D => cw_9_port, CK => N442, RN => Rst, Q 
                           => cw1_1_port, QN => net43177);
   cw1_reg_0_inst : DFFR_X1 port map( D => cw_2_port, CK => N442, RN => Rst, Q 
                           => cw1_0_port, QN => net43176);
   cw2_reg2_19_inst : DFF_X1 port map( D => n169, CK => Clk, Q => RD1_port, QN 
                           => net43175);
   cw2_reg2_18_inst : DFF_X1 port map( D => n167, CK => Clk, Q => RD2_port, QN 
                           => net43174);
   cw2_reg2_17_inst : DFF_X1 port map( D => n165, CK => Clk, Q => 
                           RegIMM_LATCH_EN_port, QN => net43173);
   cw2_reg2_16_inst : DFF_X1 port map( D => n163, CK => Clk, Q => 
                           Reg_RD1_EN_port, QN => net43172);
   cw2_reg2_15_inst : DFF_X1 port map( D => n161, CK => Clk, Q => cw2_15_port, 
                           QN => net43171);
   cw2_reg2_14_inst : DFF_X1 port map( D => n159, CK => Clk, Q => cw2_14_port, 
                           QN => net43170);
   cw2_reg2_13_inst : DFF_X1 port map( D => n157, CK => Clk, Q => cw2_13_port, 
                           QN => net43169);
   cw2_reg2_12_inst : DFF_X1 port map( D => n155, CK => Clk, Q => cw2_12_port, 
                           QN => net43168);
   cw2_reg2_11_inst : DFF_X1 port map( D => n153, CK => Clk, Q => cw2_11_port, 
                           QN => net43167);
   cw2_reg2_10_inst : DFF_X1 port map( D => n151, CK => Clk, Q => cw2_10_port, 
                           QN => net43166);
   cw2_reg2_9_inst : DFF_X1 port map( D => n149, CK => Clk, Q => cw2_9_port, QN
                           => net43165);
   cw2_reg2_8_inst : DFF_X1 port map( D => n147, CK => Clk, Q => cw2_8_port, QN
                           => net43164);
   cw2_reg2_7_inst : DFF_X1 port map( D => n145, CK => Clk, Q => cw2_7_port, QN
                           => net43163);
   cw2_reg2_6_inst : DFF_X1 port map( D => n143, CK => Clk, Q => cw2_6_port, QN
                           => net43162);
   cw2_reg2_5_inst : DFF_X1 port map( D => n141, CK => Clk, Q => cw2_5_port, QN
                           => net43161);
   cw2_reg2_4_inst : DFF_X1 port map( D => n139, CK => Clk, Q => cw2_4_port, QN
                           => net43160);
   cw2_reg2_3_inst : DFF_X1 port map( D => n137, CK => Clk, Q => cw2_3_port, QN
                           => net43159);
   cw2_reg2_2_inst : DFF_X1 port map( D => n135, CK => Clk, Q => cw2_2_port, QN
                           => net43158);
   cw2_reg2_1_inst : DFF_X1 port map( D => n133, CK => Clk, Q => cw2_1_port, QN
                           => net43157);
   cw2_reg2_0_inst : DFF_X1 port map( D => n131, CK => Clk, Q => cw2_0_port, QN
                           => net43156);
   cw1_reg2_20_inst : DFF_X1 port map( D => n129, CK => Clk, Q => 
                           IR_LATCH_EN_port, QN => net43155);
   cw1_reg2_19_inst : DFF_X1 port map( D => n127, CK => Clk, Q => cw1_19_port, 
                           QN => net43154);
   cw2_reg_19_inst : DFFR_X1 port map( D => cw1_19_port, CK => N442, RN => Rst,
                           Q => RD1_port, QN => net43153);
   cw1_reg2_18_inst : DFF_X1 port map( D => n124, CK => Clk, Q => cw1_18_port, 
                           QN => net43152);
   cw2_reg_18_inst : DFFR_X1 port map( D => cw1_18_port, CK => N442, RN => Rst,
                           Q => RD2_port, QN => net43151);
   cw1_reg2_17_inst : DFF_X1 port map( D => n121, CK => Clk, Q => cw1_17_port, 
                           QN => net43150);
   cw2_reg_17_inst : DFFR_X1 port map( D => cw1_17_port, CK => N442, RN => Rst,
                           Q => RegIMM_LATCH_EN_port, QN => net43149);
   cw1_reg2_16_inst : DFF_X1 port map( D => n118, CK => Clk, Q => cw1_16_port, 
                           QN => net43148);
   cw2_reg_16_inst : DFFR_X1 port map( D => cw1_16_port, CK => N442, RN => Rst,
                           Q => Reg_RD1_EN_port, QN => net43147);
   cw1_reg2_15_inst : DFF_X1 port map( D => n115, CK => Clk, Q => cw1_15_port, 
                           QN => net43146);
   cw2_reg_15_inst : DFFR_X1 port map( D => cw1_15_port, CK => N442, RN => Rst,
                           Q => cw2_15_port, QN => net43145);
   cw1_reg2_14_inst : DFF_X1 port map( D => n111, CK => Clk, Q => cw1_14_port, 
                           QN => net43144);
   cw2_reg_14_inst : DFFR_X1 port map( D => cw1_14_port, CK => N442, RN => Rst,
                           Q => cw2_14_port, QN => net43143);
   cw1_reg2_13_inst : DFF_X1 port map( D => n107, CK => Clk, Q => cw1_13_port, 
                           QN => net43142);
   cw1_reg2_12_inst : DFF_X1 port map( D => n103, CK => Clk, Q => cw1_12_port, 
                           QN => net43141);
   cw2_reg_12_inst : DFFR_X1 port map( D => cw1_12_port, CK => N442, RN => Rst,
                           Q => cw2_12_port, QN => net43140);
   cw3_reg_12_inst : DFFR_X1 port map( D => cw2_12_port, CK => N442, RN => Rst,
                           Q => Reg_RD2_EN, QN => n100);
   cw1_reg2_11_inst : DFF_X1 port map( D => n99, CK => Clk, Q => cw1_11_port, 
                           QN => net43139);
   cw2_reg_11_inst : DFFR_X1 port map( D => cw1_11_port, CK => N442, RN => Rst,
                           Q => cw2_11_port, QN => net43138);
   cw3_reg_11_inst : DFFR_X1 port map( D => cw2_11_port, CK => N442, RN => Rst,
                           Q => JUMP_en, QN => n96);
   cw1_reg2_10_inst : DFF_X1 port map( D => n95, CK => Clk, Q => cw1_10_port, 
                           QN => net43137);
   cw2_reg_10_inst : DFFR_X1 port map( D => cw1_10_port, CK => N442, RN => Rst,
                           Q => cw2_10_port, QN => net43136);
   cw3_reg_10_inst : DFFR_X1 port map( D => cw2_10_port, CK => N442, RN => Rst,
                           Q => cw3_10_port, QN => n92);
   cw4_reg_10_inst : DFFR_X1 port map( D => cw3_10_port, CK => N442, RN => Rst,
                           Q => DRAM_WE, QN => n91);
   cw1_reg2_9_inst : DFF_X1 port map( D => n90, CK => Clk, Q => cw1_9_port, QN 
                           => net43135);
   cw2_reg_9_inst : DFFR_X1 port map( D => cw1_9_port, CK => N442, RN => Rst, Q
                           => cw2_9_port, QN => net43134);
   cw3_reg_9_inst : DFFR_X1 port map( D => cw2_9_port, CK => N442, RN => Rst, Q
                           => cw3_9_port, QN => n87);
   cw1_reg2_8_inst : DFF_X1 port map( D => n85, CK => Clk, Q => cw1_8_port, QN 
                           => net43133);
   cw2_reg_8_inst : DFFR_X1 port map( D => cw1_8_port, CK => N442, RN => Rst, Q
                           => cw2_8_port, QN => net43132);
   cw3_reg_8_inst : DFFR_X1 port map( D => cw2_8_port, CK => N442, RN => Rst, Q
                           => cw3_8_port, QN => n82);
   cw1_reg2_7_inst : DFF_X1 port map( D => n80, CK => Clk, Q => cw1_7_port, QN 
                           => net43131);
   cw2_reg_7_inst : DFFR_X1 port map( D => cw1_7_port, CK => N442, RN => Rst, Q
                           => cw2_7_port, QN => net43130);
   cw3_reg_7_inst : DFFR_X1 port map( D => cw2_7_port, CK => N442, RN => Rst, Q
                           => cw3_7_port, QN => n77);
   cw1_reg2_6_inst : DFF_X1 port map( D => n75, CK => Clk, Q => cw1_6_port, QN 
                           => net43129);
   cw2_reg_6_inst : DFFR_X1 port map( D => cw1_6_port, CK => N442, RN => Rst, Q
                           => cw2_6_port, QN => net43128);
   cw3_reg_6_inst : DFFR_X1 port map( D => cw2_6_port, CK => N442, RN => Rst, Q
                           => cw3_6_port, QN => n72);
   cw4_reg_6_inst : DFFR_X1 port map( D => cw3_6_port, CK => N442, RN => Rst, Q
                           => PC_LATCH_EN, QN => n71);
   cw1_reg2_5_inst : DFF_X1 port map( D => n70, CK => Clk, Q => cw1_5_port, QN 
                           => net43127);
   cw2_reg_5_inst : DFFR_X1 port map( D => cw1_5_port, CK => N442, RN => Rst, Q
                           => cw2_5_port, QN => net43126);
   cw3_reg_5_inst : DFFR_X1 port map( D => cw2_5_port, CK => N442, RN => Rst, Q
                           => cw3_5_port, QN => n67);
   cw4_reg_5_inst : DFFR_X1 port map( D => cw3_5_port, CK => N442, RN => Rst, Q
                           => Reg_RD3_EN, QN => n66);
   cw1_reg2_4_inst : DFF_X1 port map( D => n65, CK => Clk, Q => cw1_4_port, QN 
                           => net43125);
   cw2_reg_4_inst : DFFR_X1 port map( D => cw1_4_port, CK => N442, RN => Rst, Q
                           => cw2_4_port, QN => net43124);
   cw3_reg_4_inst : DFFR_X1 port map( D => cw2_4_port, CK => N442, RN => Rst, Q
                           => cw3_4_port, QN => n62);
   cw4_reg_4_inst : DFFR_X1 port map( D => cw3_4_port, CK => N442, RN => Rst, Q
                           => write_stop_if_branch, QN => n61);
   cw1_reg2_3_inst : DFF_X1 port map( D => n60, CK => Clk, Q => cw1_3_port, QN 
                           => net43123);
   cw2_reg_3_inst : DFFR_X1 port map( D => cw1_3_port, CK => N442, RN => Rst, Q
                           => cw2_3_port, QN => net43122);
   cw3_reg_3_inst : DFFR_X1 port map( D => cw2_3_port, CK => N442, RN => Rst, Q
                           => cw3_3_port, QN => n57);
   cw4_reg_3_inst : DFFR_X1 port map( D => cw3_3_port, CK => N442, RN => Rst, Q
                           => cw4_3_port, QN => n56);
   cw1_reg2_2_inst : DFF_X1 port map( D => n54, CK => Clk, Q => cw1_2_port, QN 
                           => net43121);
   cw2_reg_2_inst : DFFR_X1 port map( D => cw1_2_port, CK => N442, RN => Rst, Q
                           => cw2_2_port, QN => net43120);
   cw3_reg_2_inst : DFFR_X1 port map( D => cw2_2_port, CK => N442, RN => Rst, Q
                           => cw3_2_port, QN => n51);
   cw4_reg_2_inst : DFFR_X1 port map( D => cw3_2_port, CK => N442, RN => Rst, Q
                           => cw4_2_port, QN => n50);
   cw5_reg_2_inst : DFFR_X1 port map( D => cw4_2_port, CK => N442, RN => Rst, Q
                           => RF_WE, QN => n49);
   cw1_reg2_1_inst : DFF_X1 port map( D => n48, CK => Clk, Q => cw1_1_port, QN 
                           => net43119);
   cw2_reg_1_inst : DFFR_X1 port map( D => cw1_1_port, CK => N442, RN => Rst, Q
                           => cw2_1_port, QN => net43118);
   cw3_reg_1_inst : DFFR_X1 port map( D => cw2_1_port, CK => N442, RN => Rst, Q
                           => cw3_1_port, QN => n45);
   cw4_reg_1_inst : DFFR_X1 port map( D => cw3_1_port, CK => N442, RN => Rst, Q
                           => cw4_1_port, QN => n44);
   cw5_reg_1_inst : DFFR_X1 port map( D => cw4_1_port, CK => N442, RN => Rst, Q
                           => WB_MUX_ADD_SEL, QN => n43);
   cw1_reg2_0_inst : DFF_X1 port map( D => n42, CK => Clk, Q => cw1_0_port, QN 
                           => net43117);
   cw2_reg_0_inst : DFFR_X1 port map( D => cw1_0_port, CK => N442, RN => Rst, Q
                           => cw2_0_port, QN => net43116);
   cw3_reg_0_inst : DFFR_X1 port map( D => cw2_0_port, CK => N442, RN => Rst, Q
                           => cw3_0_port, QN => n39);
   cw4_reg_0_inst : DFFR_X1 port map( D => cw3_0_port, CK => N442, RN => Rst, Q
                           => cw4_0_port, QN => n38);
   cw5_reg_0_inst : DFFR_X1 port map( D => cw4_0_port, CK => N442, RN => Rst, Q
                           => WR, QN => n37);
   cw3_reg_13_inst : DFFR_X2 port map( D => cw2_13_port, CK => N442, RN => Rst,
                           Q => ALU_OUTREG_EN, QN => n7);
   cw5_reg_3_inst : DFFR_X2 port map( D => cw4_3_port, CK => N442, RN => Rst, Q
                           => WB_MUX_SEL, QN => n6);
   cw3_reg_15_inst : DFFR_X2 port map( D => cw2_15_port, CK => N442, RN => Rst,
                           Q => MUXA_SEL, QN => n5);
   cw4_reg_7_inst : DFFR_X2 port map( D => cw3_7_port, CK => N442, RN => Rst, Q
                           => Alu_outreg2_en, QN => n4);
   cw3_reg_14_inst : DFFR_X2 port map( D => cw2_14_port, CK => N442, RN => Rst,
                           Q => MUXB_SEL, QN => n3);
   cw4_reg_8_inst : DFFR_X2 port map( D => cw3_8_port, CK => N442, RN => Rst, Q
                           => LMD_LATCH_EN, QN => n2);
   cw4_reg_9_inst : DFFR_X2 port map( D => cw3_9_port, CK => N442, RN => Rst, Q
                           => ALU_OUT2_SEL, QN => n1);
   cw2_reg_13_inst : DFFR_X1 port map( D => cw1_13_port, CK => N442, RN => Rst,
                           Q => cw2_13_port, QN => net43115);
   U3 : INV_X4 port map( A => Clk, ZN => N442);
   U4 : NAND2_X4 port map( A1 => n13, A2 => n12, ZN => RegAluOpCodeGen_EN_port)
                           ;
   U5 : INV_X2 port map( A => flush, ZN => n11);
   U6 : INV_X4 port map( A => n7, ZN => B2_LATCH_EN_port);
   U7 : INV_X1 port map( A => IR_LATCH_EN_port, ZN => n9);
   U8 : INV_X8 port map( A => n9, ZN => NPC1_LATCH_EN_port);
   U9 : AND2_X1 port map( A1 => cw1_11_port, A2 => n11, ZN => n99);
   U10 : AND2_X1 port map( A1 => cw1_10_port, A2 => n11, ZN => n95);
   U11 : AND2_X1 port map( A1 => cw1_9_port, A2 => n11, ZN => n90);
   U12 : AND2_X1 port map( A1 => cw1_8_port, A2 => n11, ZN => n85);
   U13 : AND2_X1 port map( A1 => cw1_7_port, A2 => n11, ZN => n80);
   U14 : AND2_X1 port map( A1 => cw1_6_port, A2 => n11, ZN => n75);
   U15 : AND2_X1 port map( A1 => cw1_5_port, A2 => n11, ZN => n70);
   U16 : AND2_X1 port map( A1 => cw1_4_port, A2 => n11, ZN => n65);
   U17 : AND2_X1 port map( A1 => cw1_3_port, A2 => n11, ZN => n60);
   U18 : AND2_X1 port map( A1 => cw1_2_port, A2 => n11, ZN => n54);
   U19 : AND2_X1 port map( A1 => cw1_1_port, A2 => n11, ZN => n48);
   U20 : AND2_X1 port map( A1 => cw1_0_port, A2 => n11, ZN => n42);
   U21 : AND2_X1 port map( A1 => RD1_port, A2 => n11, ZN => n169);
   U22 : AND2_X1 port map( A1 => RD2_port, A2 => n11, ZN => n167);
   U23 : NOR2_X1 port map( A1 => flush, A2 => n12, ZN => n165);
   U24 : NOR2_X1 port map( A1 => flush, A2 => n13, ZN => n163);
   U25 : AND2_X1 port map( A1 => cw2_15_port, A2 => n11, ZN => n161);
   U26 : AND2_X1 port map( A1 => cw2_14_port, A2 => n11, ZN => n159);
   U27 : AND2_X1 port map( A1 => cw2_13_port, A2 => n11, ZN => n157);
   U28 : AND2_X1 port map( A1 => cw2_12_port, A2 => n11, ZN => n155);
   U29 : AND2_X1 port map( A1 => cw2_11_port, A2 => n11, ZN => n153);
   U30 : AND2_X1 port map( A1 => cw2_10_port, A2 => n11, ZN => n151);
   U31 : AND2_X1 port map( A1 => cw2_9_port, A2 => n11, ZN => n149);
   U32 : AND2_X1 port map( A1 => cw2_8_port, A2 => n11, ZN => n147);
   U33 : AND2_X1 port map( A1 => cw2_7_port, A2 => n11, ZN => n145);
   U34 : AND2_X1 port map( A1 => cw2_6_port, A2 => n11, ZN => n143);
   U35 : AND2_X1 port map( A1 => cw2_5_port, A2 => n11, ZN => n141);
   U36 : AND2_X1 port map( A1 => cw2_4_port, A2 => n11, ZN => n139);
   U37 : AND2_X1 port map( A1 => cw2_3_port, A2 => n11, ZN => n137);
   U38 : AND2_X1 port map( A1 => cw2_2_port, A2 => n11, ZN => n135);
   U39 : AND2_X1 port map( A1 => cw2_1_port, A2 => n11, ZN => n133);
   U40 : AND2_X1 port map( A1 => cw2_0_port, A2 => n11, ZN => n131);
   U41 : AND2_X1 port map( A1 => NPC1_LATCH_EN_port, A2 => n11, ZN => n129);
   U42 : AND2_X1 port map( A1 => cw1_19_port, A2 => n11, ZN => n127);
   U43 : AND2_X1 port map( A1 => cw1_18_port, A2 => n11, ZN => n124);
   U44 : AND2_X1 port map( A1 => cw1_17_port, A2 => n11, ZN => n121);
   U45 : AND2_X1 port map( A1 => cw1_16_port, A2 => n11, ZN => n118);
   U46 : AND2_X1 port map( A1 => cw1_15_port, A2 => n11, ZN => n115);
   U47 : AND2_X1 port map( A1 => cw1_14_port, A2 => n11, ZN => n111);
   U48 : AND2_X1 port map( A1 => cw1_13_port, A2 => n11, ZN => n107);
   U49 : AND2_X1 port map( A1 => cw1_12_port, A2 => n11, ZN => n103);
   U50 : NAND2_X1 port map( A1 => n14, A2 => n15, ZN => cw_6_port);
   U51 : INV_X1 port map( A => cw_7_port, ZN => n15);
   U52 : NAND2_X1 port map( A1 => n16, A2 => n17, ZN => cw_7_port);
   U53 : NAND3_X1 port map( A1 => n18, A2 => n19, A3 => n20, ZN => n14);
   U54 : OR2_X1 port map( A1 => cw_5_port, A2 => cw_9_port, ZN => cw_2_port);
   U55 : NOR2_X1 port map( A1 => n21, A2 => n16, ZN => cw_9_port);
   U56 : INV_X1 port map( A => n17, ZN => cw_5_port);
   U57 : NAND2_X1 port map( A1 => n22, A2 => n17, ZN => cw_19_port);
   U58 : NOR2_X1 port map( A1 => n23, A2 => cw_18_port, ZN => n17);
   U59 : INV_X1 port map( A => n24, ZN => cw_18_port);
   U60 : AOI221_X1 port map( B1 => IR_IN(5), B2 => n25, C1 => n26, C2 => 
                           IR_IN(3), A => n27, ZN => n24);
   U61 : INV_X1 port map( A => n28, ZN => n27);
   U62 : OAI21_X1 port map( B1 => n25, B2 => n26, A => IR_IN(2), ZN => n28);
   U63 : NOR4_X1 port map( A1 => n29, A2 => n30, A3 => IR_IN(1), A4 => n31, ZN 
                           => n26);
   U64 : INV_X1 port map( A => IR_IN(5), ZN => n30);
   U65 : INV_X1 port map( A => IR_IN(0), ZN => n29);
   U66 : NOR3_X1 port map( A1 => IR_IN(0), A2 => IR_IN(3), A3 => n31, ZN => n25
                           );
   U67 : OR4_X1 port map( A1 => IR_IN(10), A2 => n32, A3 => n33, A4 => n34, ZN 
                           => n31);
   U68 : NAND4_X1 port map( A1 => n35, A2 => n19, A3 => n18, A4 => n36, ZN => 
                           n34);
   U69 : NOR2_X1 port map( A1 => IR_IN(9), A2 => IR_IN(8), ZN => n36);
   U70 : OR3_X1 port map( A1 => IR_IN(7), A2 => IR_IN(6), A3 => IR_IN(4), ZN =>
                           n33);
   U71 : OR2_X1 port map( A1 => n23, A2 => cw_4_port, ZN => cw_17_port);
   U72 : OAI21_X1 port map( B1 => IR_IN(29), B2 => n22, A => n16, ZN => 
                           cw_4_port);
   U73 : OR2_X1 port map( A1 => n23, A2 => cw_15_port, ZN => cw_14_port);
   U74 : INV_X1 port map( A => n16, ZN => cw_15_port);
   U75 : NAND2_X1 port map( A1 => n40, A2 => n41, ZN => n16);
   U76 : OAI211_X1 port map( C1 => n19, C2 => n22, A => n46, B => n47, ZN => 
                           n23);
   U77 : NOR2_X1 port map( A1 => cw_8_port, A2 => n52, ZN => n47);
   U78 : NOR4_X1 port map( A1 => n53, A2 => n21, A3 => IR_IN(31), A4 => 
                           IR_IN(27), ZN => n52);
   U79 : NAND2_X1 port map( A1 => IR_IN(30), A2 => IR_IN(29), ZN => n53);
   U80 : AND3_X1 port map( A1 => IR_IN(26), A2 => n40, A3 => IR_IN(31), ZN => 
                           cw_8_port);
   U81 : NOR4_X1 port map( A1 => n18, A2 => IR_IN(28), A3 => IR_IN(29), A4 => 
                           IR_IN(30), ZN => n40);
   U82 : MUX2_X1 port map( A => n55, B => n32, S => IR_IN(29), Z => n46);
   U83 : NAND3_X1 port map( A1 => n58, A2 => n41, A3 => n21, ZN => n32);
   U84 : INV_X1 port map( A => IR_IN(31), ZN => n41);
   U85 : NAND3_X1 port map( A1 => IR_IN(30), A2 => n21, A3 => n20, ZN => n55);
   U86 : INV_X1 port map( A => IR_IN(26), ZN => n21);
   U87 : NAND3_X1 port map( A1 => n18, A2 => n58, A3 => n20, ZN => n22);
   U88 : NOR2_X1 port map( A1 => n35, A2 => IR_IN(31), ZN => n20);
   U89 : INV_X1 port map( A => IR_IN(28), ZN => n35);
   U90 : INV_X1 port map( A => IR_IN(30), ZN => n58);
   U91 : INV_X1 port map( A => IR_IN(27), ZN => n18);
   U92 : INV_X1 port map( A => IR_IN(29), ZN => n19);
   U93 : INV_X1 port map( A => RegIMM_LATCH_EN_port, ZN => n12);
   U94 : INV_X1 port map( A => Reg_RD1_EN_port, ZN => n13);

end SYN_beh;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity mux21_N32_0 is

   port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (31 downto 0));

end mux21_N32_0;

architecture SYN_behavioural of mux21_N32_0 is

   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;

begin
   
   U1 : MUX2_X1 port map( A => A(9), B => B(9), S => SEL, Z => Y(9));
   U2 : MUX2_X1 port map( A => A(8), B => B(8), S => SEL, Z => Y(8));
   U3 : MUX2_X1 port map( A => A(7), B => B(7), S => SEL, Z => Y(7));
   U4 : MUX2_X1 port map( A => A(6), B => B(6), S => SEL, Z => Y(6));
   U5 : MUX2_X1 port map( A => A(5), B => B(5), S => SEL, Z => Y(5));
   U6 : MUX2_X1 port map( A => A(4), B => B(4), S => SEL, Z => Y(4));
   U7 : MUX2_X1 port map( A => A(3), B => B(3), S => SEL, Z => Y(3));
   U8 : MUX2_X1 port map( A => A(31), B => B(31), S => SEL, Z => Y(31));
   U9 : MUX2_X1 port map( A => A(30), B => B(30), S => SEL, Z => Y(30));
   U10 : MUX2_X1 port map( A => A(2), B => B(2), S => SEL, Z => Y(2));
   U11 : MUX2_X1 port map( A => A(29), B => B(29), S => SEL, Z => Y(29));
   U12 : MUX2_X1 port map( A => A(28), B => B(28), S => SEL, Z => Y(28));
   U13 : MUX2_X1 port map( A => A(27), B => B(27), S => SEL, Z => Y(27));
   U14 : MUX2_X1 port map( A => A(26), B => B(26), S => SEL, Z => Y(26));
   U15 : MUX2_X1 port map( A => A(25), B => B(25), S => SEL, Z => Y(25));
   U16 : MUX2_X1 port map( A => A(24), B => B(24), S => SEL, Z => Y(24));
   U17 : MUX2_X1 port map( A => A(23), B => B(23), S => SEL, Z => Y(23));
   U18 : MUX2_X1 port map( A => A(22), B => B(22), S => SEL, Z => Y(22));
   U19 : MUX2_X1 port map( A => A(21), B => B(21), S => SEL, Z => Y(21));
   U20 : MUX2_X1 port map( A => A(20), B => B(20), S => SEL, Z => Y(20));
   U21 : MUX2_X1 port map( A => A(1), B => B(1), S => SEL, Z => Y(1));
   U22 : MUX2_X1 port map( A => A(19), B => B(19), S => SEL, Z => Y(19));
   U23 : MUX2_X1 port map( A => A(18), B => B(18), S => SEL, Z => Y(18));
   U24 : MUX2_X1 port map( A => A(17), B => B(17), S => SEL, Z => Y(17));
   U25 : MUX2_X1 port map( A => A(16), B => B(16), S => SEL, Z => Y(16));
   U26 : MUX2_X1 port map( A => A(15), B => B(15), S => SEL, Z => Y(15));
   U27 : MUX2_X1 port map( A => A(14), B => B(14), S => SEL, Z => Y(14));
   U28 : MUX2_X1 port map( A => A(13), B => B(13), S => SEL, Z => Y(13));
   U29 : MUX2_X1 port map( A => A(12), B => B(12), S => SEL, Z => Y(12));
   U30 : MUX2_X1 port map( A => A(11), B => B(11), S => SEL, Z => Y(11));
   U31 : MUX2_X1 port map( A => A(10), B => B(10), S => SEL, Z => Y(10));
   U32 : MUX2_X1 port map( A => A(0), B => B(0), S => SEL, Z => Y(0));

end SYN_behavioural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity datapath_reg_size32 is

   port( clk, rst, flush, RF1, RF2, WF1, EN_regA, EN_regB, EN_regIMM, 
         EN_regALUOP, EN_regRD1, EN_regNPC2, S1, S2, EN_regRET, EN_regOUTALU, 
         EN_regB2, EN_regRD2, EN_regALU2, EN_regLMD, EN_regRD3, Sel_ret_alu, 
         Sel_alu_lmd, sel_31_rd : in std_logic;  NPC, IR_dp : in 
         std_logic_vector (31 downto 0);  OUT_DP : out std_logic_vector (31 
         downto 0);  comp_branch_i : out std_logic;  immediate_branch, ADD_mem,
         DIN_mem : out std_logic_vector (31 downto 0);  DOUT_mem : in 
         std_logic_vector (31 downto 0));

end datapath_reg_size32;

architecture SYN_behaviour of datapath_reg_size32 is

   component NOR3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component NAND3_X1
      port( A1, A2, A3 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component NOR4_X2
      port( A1, A2, A3, A4 : in std_logic;  ZN : out std_logic);
   end component;
   
   component CLKBUF_X3
      port( A : in std_logic;  Z : out std_logic);
   end component;
   
   component mux21_N5
      port( A, B : in std_logic_vector (4 downto 0);  SEL : in std_logic;  Y : 
            out std_logic_vector (4 downto 0));
   end component;
   
   component mux21_N32_1
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component registro_N5_1
      port( data : in std_logic_vector (4 downto 0);  enable, clock, clear : in
            std_logic;  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component registro_N32_1
      port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : 
            in std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component registro_N32_2
      port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : 
            in std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_N32_2
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component registro_N32_3
      port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : 
            in std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component registro_N5_2
      port( data : in std_logic_vector (4 downto 0);  enable, clock, clear : in
            std_logic;  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component registro_N32_4
      port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : 
            in std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component registro_N32_5
      port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : 
            in std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component AluOpCodeGen
      port( IR_opcode : in std_logic_vector (5 downto 0);  IR_func : in 
            std_logic_vector (10 downto 0);  AluOpCode : out std_logic_vector 
            (2 downto 0);  Add_Subn : out std_logic;  CompareCode : out 
            std_logic_vector (3 downto 0);  ShiftOpCode : out std_logic_vector 
            (2 downto 0));
   end component;
   
   component ALU_N32
      port( AluOpCode : in std_logic_vector (2 downto 0);  CompareOpCode : in 
            std_logic_vector (3 downto 0);  Add_subn : in std_logic;  
            ShiftOpCode : in std_logic_vector (2 downto 0);  DATA1, DATA2 : in 
            std_logic_vector (31 downto 0);  OUTALU, return_address : out 
            std_logic_vector (31 downto 0);  CompBranch : out std_logic);
   end component;
   
   component mux21_N32_3
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component mux21_N32_4
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component registro_N5_0
      port( data : in std_logic_vector (4 downto 0);  enable, clock, clear : in
            std_logic;  Q : out std_logic_vector (4 downto 0));
   end component;
   
   component registro_N17
      port( data : in std_logic_vector (16 downto 0);  enable, clock, clear : 
            in std_logic;  Q : out std_logic_vector (16 downto 0));
   end component;
   
   component registro_N32_6
      port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : 
            in std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component registro_N32_7
      port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : 
            in std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component registro_N32_8
      port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : 
            in std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component registro_N32_0
      port( data : in std_logic_vector (31 downto 0);  enable, clock, clear : 
            in std_logic;  Q : out std_logic_vector (31 downto 0));
   end component;
   
   component SIG_EXT_BITS32
      port( EXT_UNSIGNED, EXT_FOR_J : in std_logic;  S_IN : in std_logic_vector
            (31 downto 0);  S_OUT : out std_logic_vector (31 downto 0));
   end component;
   
   component register_file_NBIT32_row32
      port( CLK, RESET, ENABLE, RD1, RD2, WR : in std_logic;  ADD_WR, ADD_RD1, 
            ADD_RD2 : in std_logic_vector (4 downto 0);  DATAIN : in 
            std_logic_vector (31 downto 0);  OUT1, OUT2 : out std_logic_vector 
            (31 downto 0));
   end component;
   
   component DLL_X1
      port( D, GN : in std_logic;  Q : out std_logic);
   end component;
   
   component DLH_X1
      port( G, D : in std_logic;  Q : out std_logic);
   end component;
   
   signal X_Logic1_port, ADD_mem_31_port, ADD_mem_30_port, ADD_mem_29_port, 
      ADD_mem_28_port, ADD_mem_27_port, ADD_mem_26_port, ADD_mem_25_port, 
      ADD_mem_24_port, ADD_mem_23_port, ADD_mem_22_port, ADD_mem_21_port, 
      ADD_mem_20_port, ADD_mem_19_port, ADD_mem_18_port, ADD_mem_17_port, 
      ADD_mem_16_port, ADD_mem_15_port, ADD_mem_14_port, ADD_mem_13_port, 
      ADD_mem_12_port, ADD_mem_11_port, ADD_mem_10_port, ADD_mem_9_port, 
      ADD_mem_8_port, ADD_mem_7_port, ADD_mem_6_port, ADD_mem_5_port, 
      ADD_mem_4_port, ADD_mem_3_port, ADD_mem_2_port, ADD_mem_1_port, 
      ADD_mem_0_port, immediate_branch_31_port, immediate_branch_30_port, 
      immediate_branch_29_port, immediate_branch_28_port, 
      immediate_branch_27_port, immediate_branch_26_port, 
      immediate_branch_25_port, immediate_branch_24_port, 
      immediate_branch_23_port, immediate_branch_22_port, 
      immediate_branch_21_port, immediate_branch_20_port, 
      immediate_branch_19_port, immediate_branch_18_port, 
      immediate_branch_17_port, immediate_branch_16_port, 
      immediate_branch_15_port, immediate_branch_14_port, 
      immediate_branch_13_port, immediate_branch_12_port, 
      immediate_branch_11_port, immediate_branch_10_port, 
      immediate_branch_9_port, immediate_branch_8_port, immediate_branch_7_port
      , immediate_branch_6_port, immediate_branch_5_port, 
      immediate_branch_4_port, immediate_branch_3_port, immediate_branch_2_port
      , immediate_branch_1_port, immediate_branch_0_port, reset_pipe2, 
      add_w_rf_4_port, add_w_rf_3_port, add_w_rf_2_port, add_w_rf_1_port, 
      add_w_rf_0_port, alu2_lmd_31_port, alu2_lmd_30_port, alu2_lmd_29_port, 
      alu2_lmd_28_port, alu2_lmd_27_port, alu2_lmd_26_port, alu2_lmd_25_port, 
      alu2_lmd_24_port, alu2_lmd_23_port, alu2_lmd_22_port, alu2_lmd_21_port, 
      alu2_lmd_20_port, alu2_lmd_19_port, alu2_lmd_18_port, alu2_lmd_17_port, 
      alu2_lmd_16_port, alu2_lmd_15_port, alu2_lmd_14_port, alu2_lmd_13_port, 
      alu2_lmd_12_port, alu2_lmd_11_port, alu2_lmd_10_port, alu2_lmd_9_port, 
      alu2_lmd_8_port, alu2_lmd_7_port, alu2_lmd_6_port, alu2_lmd_5_port, 
      alu2_lmd_4_port, alu2_lmd_3_port, alu2_lmd_2_port, alu2_lmd_1_port, 
      alu2_lmd_0_port, A_31_port, A_30_port, A_29_port, A_28_port, A_27_port, 
      A_26_port, A_25_port, A_24_port, A_23_port, A_22_port, A_21_port, 
      A_20_port, A_19_port, A_18_port, A_17_port, A_16_port, A_15_port, 
      A_14_port, A_13_port, A_12_port, A_11_port, A_10_port, A_9_port, A_8_port
      , A_7_port, A_6_port, A_5_port, A_4_port, A_3_port, A_2_port, A_1_port, 
      A_0_port, B_31_port, B_30_port, B_29_port, B_28_port, B_27_port, 
      B_26_port, B_25_port, B_24_port, B_23_port, B_22_port, B_21_port, 
      B_20_port, B_19_port, B_18_port, B_17_port, B_16_port, B_15_port, 
      B_14_port, B_13_port, B_12_port, B_11_port, B_10_port, B_9_port, B_8_port
      , B_7_port, B_6_port, B_5_port, B_4_port, B_3_port, B_2_port, B_1_port, 
      B_0_port, jump_op, ext_31_port, ext_30_port, ext_29_port, ext_28_port, 
      ext_27_port, ext_26_port, ext_25_port, ext_24_port, ext_23_port, 
      ext_22_port, ext_21_port, ext_20_port, ext_19_port, ext_18_port, 
      ext_17_port, ext_16_port, ext_15_port, ext_14_port, ext_13_port, 
      ext_12_port, ext_11_port, ext_10_port, ext_9_port, ext_8_port, ext_7_port
      , ext_6_port, ext_5_port, ext_4_port, ext_3_port, ext_2_port, ext_1_port,
      ext_0_port, out_A_31_port, out_A_30_port, out_A_29_port, out_A_28_port, 
      out_A_27_port, out_A_26_port, out_A_25_port, out_A_24_port, out_A_23_port
      , out_A_22_port, out_A_21_port, out_A_20_port, out_A_19_port, 
      out_A_18_port, out_A_17_port, out_A_16_port, out_A_15_port, out_A_14_port
      , out_A_13_port, out_A_12_port, out_A_11_port, out_A_10_port, 
      out_A_9_port, out_A_8_port, out_A_7_port, out_A_6_port, out_A_5_port, 
      out_A_4_port, out_A_3_port, out_A_2_port, out_A_1_port, out_A_0_port, 
      out_b_31_port, out_b_30_port, out_b_29_port, out_b_28_port, out_b_27_port
      , out_b_26_port, out_b_25_port, out_b_24_port, out_b_23_port, 
      out_b_22_port, out_b_21_port, out_b_20_port, out_b_19_port, out_b_18_port
      , out_b_17_port, out_b_16_port, out_b_15_port, out_b_14_port, 
      out_b_13_port, out_b_12_port, out_b_11_port, out_b_10_port, out_b_9_port,
      out_b_8_port, out_b_7_port, out_b_6_port, out_b_5_port, out_b_4_port, 
      out_b_3_port, out_b_2_port, out_b_1_port, out_b_0_port, npc2_31_port, 
      npc2_30_port, npc2_29_port, npc2_28_port, npc2_27_port, npc2_26_port, 
      npc2_25_port, npc2_24_port, npc2_23_port, npc2_22_port, npc2_21_port, 
      npc2_20_port, npc2_19_port, npc2_18_port, npc2_17_port, npc2_16_port, 
      npc2_15_port, npc2_14_port, npc2_13_port, npc2_12_port, npc2_11_port, 
      npc2_10_port, npc2_9_port, npc2_8_port, npc2_7_port, npc2_6_port, 
      npc2_5_port, npc2_4_port, npc2_3_port, npc2_2_port, npc2_1_port, 
      npc2_0_port, aluopcode_reg_out_16_port, aluopcode_reg_out_15_port, 
      aluopcode_reg_out_14_port, aluopcode_reg_out_13_port, 
      aluopcode_reg_out_12_port, aluopcode_reg_out_11_port, 
      aluopcode_reg_out_10_port, aluopcode_reg_out_9_port, 
      aluopcode_reg_out_8_port, aluopcode_reg_out_7_port, 
      aluopcode_reg_out_6_port, aluopcode_reg_out_5_port, 
      aluopcode_reg_out_4_port, aluopcode_reg_out_3_port, 
      aluopcode_reg_out_2_port, aluopcode_reg_out_1_port, 
      aluopcode_reg_out_0_port, signal_rd_in_4_port, signal_rd_in_3_port, 
      signal_rd_in_2_port, signal_rd_in_1_port, signal_rd_in_0_port, N40, N47, 
      N49, N51, N53, N55, N56, out_rd1_4_port, out_rd1_3_port, out_rd1_2_port, 
      out_rd1_1_port, out_rd1_0_port, out_mux_1_31_port, out_mux_1_30_port, 
      out_mux_1_29_port, out_mux_1_28_port, out_mux_1_27_port, 
      out_mux_1_26_port, out_mux_1_25_port, out_mux_1_24_port, 
      out_mux_1_23_port, out_mux_1_22_port, out_mux_1_21_port, 
      out_mux_1_20_port, out_mux_1_19_port, out_mux_1_18_port, 
      out_mux_1_17_port, out_mux_1_16_port, out_mux_1_15_port, 
      out_mux_1_14_port, out_mux_1_13_port, out_mux_1_12_port, 
      out_mux_1_11_port, out_mux_1_10_port, out_mux_1_9_port, out_mux_1_8_port,
      out_mux_1_7_port, out_mux_1_6_port, out_mux_1_5_port, out_mux_1_4_port, 
      out_mux_1_3_port, out_mux_1_2_port, out_mux_1_1_port, out_mux_1_0_port, 
      out_mux_2_31_port, out_mux_2_30_port, out_mux_2_29_port, 
      out_mux_2_28_port, out_mux_2_27_port, out_mux_2_26_port, 
      out_mux_2_25_port, out_mux_2_24_port, out_mux_2_23_port, 
      out_mux_2_22_port, out_mux_2_21_port, out_mux_2_20_port, 
      out_mux_2_19_port, out_mux_2_18_port, out_mux_2_17_port, 
      out_mux_2_16_port, out_mux_2_15_port, out_mux_2_14_port, 
      out_mux_2_13_port, out_mux_2_12_port, out_mux_2_11_port, 
      out_mux_2_10_port, out_mux_2_9_port, out_mux_2_8_port, out_mux_2_7_port, 
      out_mux_2_6_port, out_mux_2_5_port, out_mux_2_4_port, out_mux_2_3_port, 
      out_mux_2_2_port, out_mux_2_1_port, out_mux_2_0_port, aluopcode_i_2_port,
      aluopcode_i_1_port, aluopcode_i_0_port, compare_code_i_3_port, 
      compare_code_i_2_port, compare_code_i_1_port, compare_code_i_0_port, 
      add_sub_i, shiftopcode_i_2_port, shiftopcode_i_1_port, 
      shiftopcode_i_0_port, reg_alu_in_31_port, reg_alu_in_30_port, 
      reg_alu_in_29_port, reg_alu_in_28_port, reg_alu_in_27_port, 
      reg_alu_in_26_port, reg_alu_in_25_port, reg_alu_in_24_port, 
      reg_alu_in_23_port, reg_alu_in_22_port, reg_alu_in_21_port, 
      reg_alu_in_20_port, reg_alu_in_19_port, reg_alu_in_18_port, 
      reg_alu_in_17_port, reg_alu_in_16_port, reg_alu_in_15_port, 
      reg_alu_in_14_port, reg_alu_in_13_port, reg_alu_in_12_port, 
      reg_alu_in_11_port, reg_alu_in_10_port, reg_alu_in_9_port, 
      reg_alu_in_8_port, reg_alu_in_7_port, reg_alu_in_6_port, 
      reg_alu_in_5_port, reg_alu_in_4_port, reg_alu_in_3_port, 
      reg_alu_in_2_port, reg_alu_in_1_port, reg_alu_in_0_port, 
      return_alu_31_port, return_alu_30_port, return_alu_29_port, 
      return_alu_28_port, return_alu_27_port, return_alu_26_port, 
      return_alu_25_port, return_alu_24_port, return_alu_23_port, 
      return_alu_22_port, return_alu_21_port, return_alu_20_port, 
      return_alu_19_port, return_alu_18_port, return_alu_17_port, 
      return_alu_16_port, return_alu_15_port, return_alu_14_port, 
      return_alu_13_port, return_alu_12_port, return_alu_11_port, 
      return_alu_10_port, return_alu_9_port, return_alu_8_port, 
      return_alu_7_port, return_alu_6_port, return_alu_5_port, 
      return_alu_4_port, return_alu_3_port, return_alu_2_port, 
      return_alu_1_port, return_alu_0_port, out_rd2_4_port, out_rd2_3_port, 
      out_rd2_2_port, out_rd2_1_port, out_rd2_0_port, return_out_31_port, 
      return_out_30_port, return_out_29_port, return_out_28_port, 
      return_out_27_port, return_out_26_port, return_out_25_port, 
      return_out_24_port, return_out_23_port, return_out_22_port, 
      return_out_21_port, return_out_20_port, return_out_19_port, 
      return_out_18_port, return_out_17_port, return_out_16_port, 
      return_out_15_port, return_out_14_port, return_out_13_port, 
      return_out_12_port, return_out_11_port, return_out_10_port, 
      return_out_9_port, return_out_8_port, return_out_7_port, 
      return_out_6_port, return_out_5_port, return_out_4_port, 
      return_out_3_port, return_out_2_port, return_out_1_port, 
      return_out_0_port, out_ret_alu_31_port, out_ret_alu_30_port, 
      out_ret_alu_29_port, out_ret_alu_28_port, out_ret_alu_27_port, 
      out_ret_alu_26_port, out_ret_alu_25_port, out_ret_alu_24_port, 
      out_ret_alu_23_port, out_ret_alu_22_port, out_ret_alu_21_port, 
      out_ret_alu_20_port, out_ret_alu_19_port, out_ret_alu_18_port, 
      out_ret_alu_17_port, out_ret_alu_16_port, out_ret_alu_15_port, 
      out_ret_alu_14_port, out_ret_alu_13_port, out_ret_alu_12_port, 
      out_ret_alu_11_port, out_ret_alu_10_port, out_ret_alu_9_port, 
      out_ret_alu_8_port, out_ret_alu_7_port, out_ret_alu_6_port, 
      out_ret_alu_5_port, out_ret_alu_4_port, out_ret_alu_3_port, 
      out_ret_alu_2_port, out_ret_alu_1_port, out_ret_alu_0_port, alu2_31_port,
      alu2_30_port, alu2_29_port, alu2_28_port, alu2_27_port, alu2_26_port, 
      alu2_25_port, alu2_24_port, alu2_23_port, alu2_22_port, alu2_21_port, 
      alu2_20_port, alu2_19_port, alu2_18_port, alu2_17_port, alu2_16_port, 
      alu2_15_port, alu2_14_port, alu2_13_port, alu2_12_port, alu2_11_port, 
      alu2_10_port, alu2_9_port, alu2_8_port, alu2_7_port, alu2_6_port, 
      alu2_5_port, alu2_4_port, alu2_3_port, alu2_2_port, alu2_1_port, 
      alu2_0_port, lmd_31_port, lmd_30_port, lmd_29_port, lmd_28_port, 
      lmd_27_port, lmd_26_port, lmd_25_port, lmd_24_port, lmd_23_port, 
      lmd_22_port, lmd_21_port, lmd_20_port, lmd_19_port, lmd_18_port, 
      lmd_17_port, lmd_16_port, lmd_15_port, lmd_14_port, lmd_13_port, 
      lmd_12_port, lmd_11_port, lmd_10_port, lmd_9_port, lmd_8_port, lmd_7_port
      , lmd_6_port, lmd_5_port, lmd_4_port, lmd_3_port, lmd_2_port, lmd_1_port,
      lmd_0_port, rd3_4_port, rd3_3_port, rd3_2_port, rd3_1_port, rd3_0_port, 
      n1, n2, n3, n4, n5, n6, n7, n8 : std_logic;

begin
   OUT_DP <= ( ADD_mem_31_port, ADD_mem_30_port, ADD_mem_29_port, 
      ADD_mem_28_port, ADD_mem_27_port, ADD_mem_26_port, ADD_mem_25_port, 
      ADD_mem_24_port, ADD_mem_23_port, ADD_mem_22_port, ADD_mem_21_port, 
      ADD_mem_20_port, ADD_mem_19_port, ADD_mem_18_port, ADD_mem_17_port, 
      ADD_mem_16_port, ADD_mem_15_port, ADD_mem_14_port, ADD_mem_13_port, 
      ADD_mem_12_port, ADD_mem_11_port, ADD_mem_10_port, ADD_mem_9_port, 
      ADD_mem_8_port, ADD_mem_7_port, ADD_mem_6_port, ADD_mem_5_port, 
      ADD_mem_4_port, ADD_mem_3_port, ADD_mem_2_port, ADD_mem_1_port, 
      ADD_mem_0_port );
   immediate_branch <= ( immediate_branch_31_port, immediate_branch_30_port, 
      immediate_branch_29_port, immediate_branch_28_port, 
      immediate_branch_27_port, immediate_branch_26_port, 
      immediate_branch_25_port, immediate_branch_24_port, 
      immediate_branch_23_port, immediate_branch_22_port, 
      immediate_branch_21_port, immediate_branch_20_port, 
      immediate_branch_19_port, immediate_branch_18_port, 
      immediate_branch_17_port, immediate_branch_16_port, 
      immediate_branch_15_port, immediate_branch_14_port, 
      immediate_branch_13_port, immediate_branch_12_port, 
      immediate_branch_11_port, immediate_branch_10_port, 
      immediate_branch_9_port, immediate_branch_8_port, immediate_branch_7_port
      , immediate_branch_6_port, immediate_branch_5_port, 
      immediate_branch_4_port, immediate_branch_3_port, immediate_branch_2_port
      , immediate_branch_1_port, immediate_branch_0_port );
   ADD_mem <= ( ADD_mem_31_port, ADD_mem_30_port, ADD_mem_29_port, 
      ADD_mem_28_port, ADD_mem_27_port, ADD_mem_26_port, ADD_mem_25_port, 
      ADD_mem_24_port, ADD_mem_23_port, ADD_mem_22_port, ADD_mem_21_port, 
      ADD_mem_20_port, ADD_mem_19_port, ADD_mem_18_port, ADD_mem_17_port, 
      ADD_mem_16_port, ADD_mem_15_port, ADD_mem_14_port, ADD_mem_13_port, 
      ADD_mem_12_port, ADD_mem_11_port, ADD_mem_10_port, ADD_mem_9_port, 
      ADD_mem_8_port, ADD_mem_7_port, ADD_mem_6_port, ADD_mem_5_port, 
      ADD_mem_4_port, ADD_mem_3_port, ADD_mem_2_port, ADD_mem_1_port, 
      ADD_mem_0_port );
   
   X_Logic1_port <= '1';
   jump_op_reg : DLH_X1 port map( G => N56, D => N40, Q => jump_op);
   signal_rd_in_reg_4_inst : DLL_X1 port map( D => N55, GN => N56, Q => 
                           signal_rd_in_4_port);
   signal_rd_in_reg_3_inst : DLL_X1 port map( D => N53, GN => N56, Q => 
                           signal_rd_in_3_port);
   signal_rd_in_reg_2_inst : DLL_X1 port map( D => N51, GN => N56, Q => 
                           signal_rd_in_2_port);
   signal_rd_in_reg_1_inst : DLL_X1 port map( D => N49, GN => N56, Q => 
                           signal_rd_in_1_port);
   signal_rd_in_reg_0_inst : DLL_X1 port map( D => N47, GN => N56, Q => 
                           signal_rd_in_0_port);
   rf : register_file_NBIT32_row32 port map( CLK => clk, RESET => rst, ENABLE 
                           => X_Logic1_port, RD1 => RF1, RD2 => RF2, WR => WF1,
                           ADD_WR(4) => add_w_rf_4_port, ADD_WR(3) => 
                           add_w_rf_3_port, ADD_WR(2) => add_w_rf_2_port, 
                           ADD_WR(1) => add_w_rf_1_port, ADD_WR(0) => 
                           add_w_rf_0_port, ADD_RD1(4) => IR_dp(25), ADD_RD1(3)
                           => IR_dp(24), ADD_RD1(2) => IR_dp(23), ADD_RD1(1) =>
                           IR_dp(22), ADD_RD1(0) => IR_dp(21), ADD_RD2(4) => 
                           IR_dp(20), ADD_RD2(3) => IR_dp(19), ADD_RD2(2) => 
                           IR_dp(18), ADD_RD2(1) => IR_dp(17), ADD_RD2(0) => 
                           IR_dp(16), DATAIN(31) => alu2_lmd_31_port, 
                           DATAIN(30) => alu2_lmd_30_port, DATAIN(29) => 
                           alu2_lmd_29_port, DATAIN(28) => alu2_lmd_28_port, 
                           DATAIN(27) => alu2_lmd_27_port, DATAIN(26) => 
                           alu2_lmd_26_port, DATAIN(25) => alu2_lmd_25_port, 
                           DATAIN(24) => alu2_lmd_24_port, DATAIN(23) => 
                           alu2_lmd_23_port, DATAIN(22) => alu2_lmd_22_port, 
                           DATAIN(21) => alu2_lmd_21_port, DATAIN(20) => 
                           alu2_lmd_20_port, DATAIN(19) => alu2_lmd_19_port, 
                           DATAIN(18) => alu2_lmd_18_port, DATAIN(17) => 
                           alu2_lmd_17_port, DATAIN(16) => alu2_lmd_16_port, 
                           DATAIN(15) => alu2_lmd_15_port, DATAIN(14) => 
                           alu2_lmd_14_port, DATAIN(13) => alu2_lmd_13_port, 
                           DATAIN(12) => alu2_lmd_12_port, DATAIN(11) => 
                           alu2_lmd_11_port, DATAIN(10) => alu2_lmd_10_port, 
                           DATAIN(9) => alu2_lmd_9_port, DATAIN(8) => 
                           alu2_lmd_8_port, DATAIN(7) => alu2_lmd_7_port, 
                           DATAIN(6) => alu2_lmd_6_port, DATAIN(5) => 
                           alu2_lmd_5_port, DATAIN(4) => alu2_lmd_4_port, 
                           DATAIN(3) => alu2_lmd_3_port, DATAIN(2) => 
                           alu2_lmd_2_port, DATAIN(1) => alu2_lmd_1_port, 
                           DATAIN(0) => alu2_lmd_0_port, OUT1(31) => A_31_port,
                           OUT1(30) => A_30_port, OUT1(29) => A_29_port, 
                           OUT1(28) => A_28_port, OUT1(27) => A_27_port, 
                           OUT1(26) => A_26_port, OUT1(25) => A_25_port, 
                           OUT1(24) => A_24_port, OUT1(23) => A_23_port, 
                           OUT1(22) => A_22_port, OUT1(21) => A_21_port, 
                           OUT1(20) => A_20_port, OUT1(19) => A_19_port, 
                           OUT1(18) => A_18_port, OUT1(17) => A_17_port, 
                           OUT1(16) => A_16_port, OUT1(15) => A_15_port, 
                           OUT1(14) => A_14_port, OUT1(13) => A_13_port, 
                           OUT1(12) => A_12_port, OUT1(11) => A_11_port, 
                           OUT1(10) => A_10_port, OUT1(9) => A_9_port, OUT1(8) 
                           => A_8_port, OUT1(7) => A_7_port, OUT1(6) => 
                           A_6_port, OUT1(5) => A_5_port, OUT1(4) => A_4_port, 
                           OUT1(3) => A_3_port, OUT1(2) => A_2_port, OUT1(1) =>
                           A_1_port, OUT1(0) => A_0_port, OUT2(31) => B_31_port
                           , OUT2(30) => B_30_port, OUT2(29) => B_29_port, 
                           OUT2(28) => B_28_port, OUT2(27) => B_27_port, 
                           OUT2(26) => B_26_port, OUT2(25) => B_25_port, 
                           OUT2(24) => B_24_port, OUT2(23) => B_23_port, 
                           OUT2(22) => B_22_port, OUT2(21) => B_21_port, 
                           OUT2(20) => B_20_port, OUT2(19) => B_19_port, 
                           OUT2(18) => B_18_port, OUT2(17) => B_17_port, 
                           OUT2(16) => B_16_port, OUT2(15) => B_15_port, 
                           OUT2(14) => B_14_port, OUT2(13) => B_13_port, 
                           OUT2(12) => B_12_port, OUT2(11) => B_11_port, 
                           OUT2(10) => B_10_port, OUT2(9) => B_9_port, OUT2(8) 
                           => B_8_port, OUT2(7) => B_7_port, OUT2(6) => 
                           B_6_port, OUT2(5) => B_5_port, OUT2(4) => B_4_port, 
                           OUT2(3) => B_3_port, OUT2(2) => B_2_port, OUT2(1) =>
                           B_1_port, OUT2(0) => B_0_port);
   estensione_segno : SIG_EXT_BITS32 port map( EXT_UNSIGNED => X_Logic1_port, 
                           EXT_FOR_J => jump_op, S_IN(31) => IR_dp(31), 
                           S_IN(30) => IR_dp(30), S_IN(29) => IR_dp(29), 
                           S_IN(28) => IR_dp(28), S_IN(27) => IR_dp(27), 
                           S_IN(26) => IR_dp(26), S_IN(25) => IR_dp(25), 
                           S_IN(24) => IR_dp(24), S_IN(23) => IR_dp(23), 
                           S_IN(22) => IR_dp(22), S_IN(21) => IR_dp(21), 
                           S_IN(20) => IR_dp(20), S_IN(19) => IR_dp(19), 
                           S_IN(18) => IR_dp(18), S_IN(17) => IR_dp(17), 
                           S_IN(16) => IR_dp(16), S_IN(15) => IR_dp(15), 
                           S_IN(14) => IR_dp(14), S_IN(13) => IR_dp(13), 
                           S_IN(12) => IR_dp(12), S_IN(11) => IR_dp(11), 
                           S_IN(10) => IR_dp(10), S_IN(9) => IR_dp(9), S_IN(8) 
                           => IR_dp(8), S_IN(7) => IR_dp(7), S_IN(6) => 
                           IR_dp(6), S_IN(5) => IR_dp(5), S_IN(4) => IR_dp(4), 
                           S_IN(3) => IR_dp(3), S_IN(2) => IR_dp(2), S_IN(1) =>
                           IR_dp(1), S_IN(0) => IR_dp(0), S_OUT(31) => 
                           ext_31_port, S_OUT(30) => ext_30_port, S_OUT(29) => 
                           ext_29_port, S_OUT(28) => ext_28_port, S_OUT(27) => 
                           ext_27_port, S_OUT(26) => ext_26_port, S_OUT(25) => 
                           ext_25_port, S_OUT(24) => ext_24_port, S_OUT(23) => 
                           ext_23_port, S_OUT(22) => ext_22_port, S_OUT(21) => 
                           ext_21_port, S_OUT(20) => ext_20_port, S_OUT(19) => 
                           ext_19_port, S_OUT(18) => ext_18_port, S_OUT(17) => 
                           ext_17_port, S_OUT(16) => ext_16_port, S_OUT(15) => 
                           ext_15_port, S_OUT(14) => ext_14_port, S_OUT(13) => 
                           ext_13_port, S_OUT(12) => ext_12_port, S_OUT(11) => 
                           ext_11_port, S_OUT(10) => ext_10_port, S_OUT(9) => 
                           ext_9_port, S_OUT(8) => ext_8_port, S_OUT(7) => 
                           ext_7_port, S_OUT(6) => ext_6_port, S_OUT(5) => 
                           ext_5_port, S_OUT(4) => ext_4_port, S_OUT(3) => 
                           ext_3_port, S_OUT(2) => ext_2_port, S_OUT(1) => 
                           ext_1_port, S_OUT(0) => ext_0_port);
   reg_A : registro_N32_0 port map( data(31) => A_31_port, data(30) => 
                           A_30_port, data(29) => A_29_port, data(28) => 
                           A_28_port, data(27) => A_27_port, data(26) => 
                           A_26_port, data(25) => A_25_port, data(24) => 
                           A_24_port, data(23) => A_23_port, data(22) => 
                           A_22_port, data(21) => A_21_port, data(20) => 
                           A_20_port, data(19) => A_19_port, data(18) => 
                           A_18_port, data(17) => A_17_port, data(16) => 
                           A_16_port, data(15) => A_15_port, data(14) => 
                           A_14_port, data(13) => A_13_port, data(12) => 
                           A_12_port, data(11) => A_11_port, data(10) => 
                           A_10_port, data(9) => A_9_port, data(8) => A_8_port,
                           data(7) => A_7_port, data(6) => A_6_port, data(5) =>
                           A_5_port, data(4) => A_4_port, data(3) => A_3_port, 
                           data(2) => A_2_port, data(1) => A_1_port, data(0) =>
                           A_0_port, enable => EN_regA, clock => clk, clear => 
                           n1, Q(31) => out_A_31_port, Q(30) => out_A_30_port, 
                           Q(29) => out_A_29_port, Q(28) => out_A_28_port, 
                           Q(27) => out_A_27_port, Q(26) => out_A_26_port, 
                           Q(25) => out_A_25_port, Q(24) => out_A_24_port, 
                           Q(23) => out_A_23_port, Q(22) => out_A_22_port, 
                           Q(21) => out_A_21_port, Q(20) => out_A_20_port, 
                           Q(19) => out_A_19_port, Q(18) => out_A_18_port, 
                           Q(17) => out_A_17_port, Q(16) => out_A_16_port, 
                           Q(15) => out_A_15_port, Q(14) => out_A_14_port, 
                           Q(13) => out_A_13_port, Q(12) => out_A_12_port, 
                           Q(11) => out_A_11_port, Q(10) => out_A_10_port, Q(9)
                           => out_A_9_port, Q(8) => out_A_8_port, Q(7) => 
                           out_A_7_port, Q(6) => out_A_6_port, Q(5) => 
                           out_A_5_port, Q(4) => out_A_4_port, Q(3) => 
                           out_A_3_port, Q(2) => out_A_2_port, Q(1) => 
                           out_A_1_port, Q(0) => out_A_0_port);
   reg_B : registro_N32_8 port map( data(31) => B_31_port, data(30) => 
                           B_30_port, data(29) => B_29_port, data(28) => 
                           B_28_port, data(27) => B_27_port, data(26) => 
                           B_26_port, data(25) => B_25_port, data(24) => 
                           B_24_port, data(23) => B_23_port, data(22) => 
                           B_22_port, data(21) => B_21_port, data(20) => 
                           B_20_port, data(19) => B_19_port, data(18) => 
                           B_18_port, data(17) => B_17_port, data(16) => 
                           B_16_port, data(15) => B_15_port, data(14) => 
                           B_14_port, data(13) => B_13_port, data(12) => 
                           B_12_port, data(11) => B_11_port, data(10) => 
                           B_10_port, data(9) => B_9_port, data(8) => B_8_port,
                           data(7) => B_7_port, data(6) => B_6_port, data(5) =>
                           B_5_port, data(4) => B_4_port, data(3) => B_3_port, 
                           data(2) => B_2_port, data(1) => B_1_port, data(0) =>
                           B_0_port, enable => EN_regB, clock => clk, clear => 
                           n1, Q(31) => out_b_31_port, Q(30) => out_b_30_port, 
                           Q(29) => out_b_29_port, Q(28) => out_b_28_port, 
                           Q(27) => out_b_27_port, Q(26) => out_b_26_port, 
                           Q(25) => out_b_25_port, Q(24) => out_b_24_port, 
                           Q(23) => out_b_23_port, Q(22) => out_b_22_port, 
                           Q(21) => out_b_21_port, Q(20) => out_b_20_port, 
                           Q(19) => out_b_19_port, Q(18) => out_b_18_port, 
                           Q(17) => out_b_17_port, Q(16) => out_b_16_port, 
                           Q(15) => out_b_15_port, Q(14) => out_b_14_port, 
                           Q(13) => out_b_13_port, Q(12) => out_b_12_port, 
                           Q(11) => out_b_11_port, Q(10) => out_b_10_port, Q(9)
                           => out_b_9_port, Q(8) => out_b_8_port, Q(7) => 
                           out_b_7_port, Q(6) => out_b_6_port, Q(5) => 
                           out_b_5_port, Q(4) => out_b_4_port, Q(3) => 
                           out_b_3_port, Q(2) => out_b_2_port, Q(1) => 
                           out_b_1_port, Q(0) => out_b_0_port);
   reg_NPC2 : registro_N32_7 port map( data(31) => NPC(31), data(30) => NPC(30)
                           , data(29) => NPC(29), data(28) => NPC(28), data(27)
                           => NPC(27), data(26) => NPC(26), data(25) => NPC(25)
                           , data(24) => NPC(24), data(23) => NPC(23), data(22)
                           => NPC(22), data(21) => NPC(21), data(20) => NPC(20)
                           , data(19) => NPC(19), data(18) => NPC(18), data(17)
                           => NPC(17), data(16) => NPC(16), data(15) => NPC(15)
                           , data(14) => NPC(14), data(13) => NPC(13), data(12)
                           => NPC(12), data(11) => NPC(11), data(10) => NPC(10)
                           , data(9) => NPC(9), data(8) => NPC(8), data(7) => 
                           NPC(7), data(6) => NPC(6), data(5) => NPC(5), 
                           data(4) => NPC(4), data(3) => NPC(3), data(2) => 
                           NPC(2), data(1) => NPC(1), data(0) => NPC(0), enable
                           => EN_regNPC2, clock => clk, clear => rst, Q(31) => 
                           npc2_31_port, Q(30) => npc2_30_port, Q(29) => 
                           npc2_29_port, Q(28) => npc2_28_port, Q(27) => 
                           npc2_27_port, Q(26) => npc2_26_port, Q(25) => 
                           npc2_25_port, Q(24) => npc2_24_port, Q(23) => 
                           npc2_23_port, Q(22) => npc2_22_port, Q(21) => 
                           npc2_21_port, Q(20) => npc2_20_port, Q(19) => 
                           npc2_19_port, Q(18) => npc2_18_port, Q(17) => 
                           npc2_17_port, Q(16) => npc2_16_port, Q(15) => 
                           npc2_15_port, Q(14) => npc2_14_port, Q(13) => 
                           npc2_13_port, Q(12) => npc2_12_port, Q(11) => 
                           npc2_11_port, Q(10) => npc2_10_port, Q(9) => 
                           npc2_9_port, Q(8) => npc2_8_port, Q(7) => 
                           npc2_7_port, Q(6) => npc2_6_port, Q(5) => 
                           npc2_5_port, Q(4) => npc2_4_port, Q(3) => 
                           npc2_3_port, Q(2) => npc2_2_port, Q(1) => 
                           npc2_1_port, Q(0) => npc2_0_port);
   reg_IMMEDIATE : registro_N32_6 port map( data(31) => ext_31_port, data(30) 
                           => ext_30_port, data(29) => ext_29_port, data(28) =>
                           ext_28_port, data(27) => ext_27_port, data(26) => 
                           ext_26_port, data(25) => ext_25_port, data(24) => 
                           ext_24_port, data(23) => ext_23_port, data(22) => 
                           ext_22_port, data(21) => ext_21_port, data(20) => 
                           ext_20_port, data(19) => ext_19_port, data(18) => 
                           ext_18_port, data(17) => ext_17_port, data(16) => 
                           ext_16_port, data(15) => ext_15_port, data(14) => 
                           ext_14_port, data(13) => ext_13_port, data(12) => 
                           ext_12_port, data(11) => ext_11_port, data(10) => 
                           ext_10_port, data(9) => ext_9_port, data(8) => 
                           ext_8_port, data(7) => ext_7_port, data(6) => 
                           ext_6_port, data(5) => ext_5_port, data(4) => 
                           ext_4_port, data(3) => ext_3_port, data(2) => 
                           ext_2_port, data(1) => ext_1_port, data(0) => 
                           ext_0_port, enable => EN_regIMM, clock => clk, clear
                           => rst, Q(31) => immediate_branch_31_port, Q(30) => 
                           immediate_branch_30_port, Q(29) => 
                           immediate_branch_29_port, Q(28) => 
                           immediate_branch_28_port, Q(27) => 
                           immediate_branch_27_port, Q(26) => 
                           immediate_branch_26_port, Q(25) => 
                           immediate_branch_25_port, Q(24) => 
                           immediate_branch_24_port, Q(23) => 
                           immediate_branch_23_port, Q(22) => 
                           immediate_branch_22_port, Q(21) => 
                           immediate_branch_21_port, Q(20) => 
                           immediate_branch_20_port, Q(19) => 
                           immediate_branch_19_port, Q(18) => 
                           immediate_branch_18_port, Q(17) => 
                           immediate_branch_17_port, Q(16) => 
                           immediate_branch_16_port, Q(15) => 
                           immediate_branch_15_port, Q(14) => 
                           immediate_branch_14_port, Q(13) => 
                           immediate_branch_13_port, Q(12) => 
                           immediate_branch_12_port, Q(11) => 
                           immediate_branch_11_port, Q(10) => 
                           immediate_branch_10_port, Q(9) => 
                           immediate_branch_9_port, Q(8) => 
                           immediate_branch_8_port, Q(7) => 
                           immediate_branch_7_port, Q(6) => 
                           immediate_branch_6_port, Q(5) => 
                           immediate_branch_5_port, Q(4) => 
                           immediate_branch_4_port, Q(3) => 
                           immediate_branch_3_port, Q(2) => 
                           immediate_branch_2_port, Q(1) => 
                           immediate_branch_1_port, Q(0) => 
                           immediate_branch_0_port);
   reg_aluopcode : registro_N17 port map( data(16) => IR_dp(31), data(15) => 
                           IR_dp(30), data(14) => IR_dp(29), data(13) => 
                           IR_dp(28), data(12) => IR_dp(27), data(11) => 
                           IR_dp(26), data(10) => IR_dp(10), data(9) => 
                           IR_dp(9), data(8) => IR_dp(8), data(7) => IR_dp(7), 
                           data(6) => IR_dp(6), data(5) => IR_dp(5), data(4) =>
                           IR_dp(4), data(3) => IR_dp(3), data(2) => IR_dp(2), 
                           data(1) => IR_dp(1), data(0) => IR_dp(0), enable => 
                           EN_regALUOP, clock => clk, clear => rst, Q(16) => 
                           aluopcode_reg_out_16_port, Q(15) => 
                           aluopcode_reg_out_15_port, Q(14) => 
                           aluopcode_reg_out_14_port, Q(13) => 
                           aluopcode_reg_out_13_port, Q(12) => 
                           aluopcode_reg_out_12_port, Q(11) => 
                           aluopcode_reg_out_11_port, Q(10) => 
                           aluopcode_reg_out_10_port, Q(9) => 
                           aluopcode_reg_out_9_port, Q(8) => 
                           aluopcode_reg_out_8_port, Q(7) => 
                           aluopcode_reg_out_7_port, Q(6) => 
                           aluopcode_reg_out_6_port, Q(5) => 
                           aluopcode_reg_out_5_port, Q(4) => 
                           aluopcode_reg_out_4_port, Q(3) => 
                           aluopcode_reg_out_3_port, Q(2) => 
                           aluopcode_reg_out_2_port, Q(1) => 
                           aluopcode_reg_out_1_port, Q(0) => 
                           aluopcode_reg_out_0_port);
   reg_rd1 : registro_N5_0 port map( data(4) => signal_rd_in_4_port, data(3) =>
                           signal_rd_in_3_port, data(2) => signal_rd_in_2_port,
                           data(1) => signal_rd_in_1_port, data(0) => 
                           signal_rd_in_0_port, enable => EN_regRD1, clock => 
                           clk, clear => n1, Q(4) => out_rd1_4_port, Q(3) => 
                           out_rd1_3_port, Q(2) => out_rd1_2_port, Q(1) => 
                           out_rd1_1_port, Q(0) => out_rd1_0_port);
   mux_in1_A : mux21_N32_4 port map( A(31) => out_A_31_port, A(30) => 
                           out_A_30_port, A(29) => out_A_29_port, A(28) => 
                           out_A_28_port, A(27) => out_A_27_port, A(26) => 
                           out_A_26_port, A(25) => out_A_25_port, A(24) => 
                           out_A_24_port, A(23) => out_A_23_port, A(22) => 
                           out_A_22_port, A(21) => out_A_21_port, A(20) => 
                           out_A_20_port, A(19) => out_A_19_port, A(18) => 
                           out_A_18_port, A(17) => out_A_17_port, A(16) => 
                           out_A_16_port, A(15) => out_A_15_port, A(14) => 
                           out_A_14_port, A(13) => out_A_13_port, A(12) => 
                           out_A_12_port, A(11) => out_A_11_port, A(10) => 
                           out_A_10_port, A(9) => out_A_9_port, A(8) => 
                           out_A_8_port, A(7) => out_A_7_port, A(6) => 
                           out_A_6_port, A(5) => out_A_5_port, A(4) => 
                           out_A_4_port, A(3) => out_A_3_port, A(2) => 
                           out_A_2_port, A(1) => out_A_1_port, A(0) => 
                           out_A_0_port, B(31) => npc2_31_port, B(30) => 
                           npc2_30_port, B(29) => npc2_29_port, B(28) => 
                           npc2_28_port, B(27) => npc2_27_port, B(26) => 
                           npc2_26_port, B(25) => npc2_25_port, B(24) => 
                           npc2_24_port, B(23) => npc2_23_port, B(22) => 
                           npc2_22_port, B(21) => npc2_21_port, B(20) => 
                           npc2_20_port, B(19) => npc2_19_port, B(18) => 
                           npc2_18_port, B(17) => npc2_17_port, B(16) => 
                           npc2_16_port, B(15) => npc2_15_port, B(14) => 
                           npc2_14_port, B(13) => npc2_13_port, B(12) => 
                           npc2_12_port, B(11) => npc2_11_port, B(10) => 
                           npc2_10_port, B(9) => npc2_9_port, B(8) => 
                           npc2_8_port, B(7) => npc2_7_port, B(6) => 
                           npc2_6_port, B(5) => npc2_5_port, B(4) => 
                           npc2_4_port, B(3) => npc2_3_port, B(2) => 
                           npc2_2_port, B(1) => npc2_1_port, B(0) => 
                           npc2_0_port, SEL => S1, Y(31) => out_mux_1_31_port, 
                           Y(30) => out_mux_1_30_port, Y(29) => 
                           out_mux_1_29_port, Y(28) => out_mux_1_28_port, Y(27)
                           => out_mux_1_27_port, Y(26) => out_mux_1_26_port, 
                           Y(25) => out_mux_1_25_port, Y(24) => 
                           out_mux_1_24_port, Y(23) => out_mux_1_23_port, Y(22)
                           => out_mux_1_22_port, Y(21) => out_mux_1_21_port, 
                           Y(20) => out_mux_1_20_port, Y(19) => 
                           out_mux_1_19_port, Y(18) => out_mux_1_18_port, Y(17)
                           => out_mux_1_17_port, Y(16) => out_mux_1_16_port, 
                           Y(15) => out_mux_1_15_port, Y(14) => 
                           out_mux_1_14_port, Y(13) => out_mux_1_13_port, Y(12)
                           => out_mux_1_12_port, Y(11) => out_mux_1_11_port, 
                           Y(10) => out_mux_1_10_port, Y(9) => out_mux_1_9_port
                           , Y(8) => out_mux_1_8_port, Y(7) => out_mux_1_7_port
                           , Y(6) => out_mux_1_6_port, Y(5) => out_mux_1_5_port
                           , Y(4) => out_mux_1_4_port, Y(3) => out_mux_1_3_port
                           , Y(2) => out_mux_1_2_port, Y(1) => out_mux_1_1_port
                           , Y(0) => out_mux_1_0_port);
   mux_in1_B : mux21_N32_3 port map( A(31) => out_b_31_port, A(30) => 
                           out_b_30_port, A(29) => out_b_29_port, A(28) => 
                           out_b_28_port, A(27) => out_b_27_port, A(26) => 
                           out_b_26_port, A(25) => out_b_25_port, A(24) => 
                           out_b_24_port, A(23) => out_b_23_port, A(22) => 
                           out_b_22_port, A(21) => out_b_21_port, A(20) => 
                           out_b_20_port, A(19) => out_b_19_port, A(18) => 
                           out_b_18_port, A(17) => out_b_17_port, A(16) => 
                           out_b_16_port, A(15) => out_b_15_port, A(14) => 
                           out_b_14_port, A(13) => out_b_13_port, A(12) => 
                           out_b_12_port, A(11) => out_b_11_port, A(10) => 
                           out_b_10_port, A(9) => out_b_9_port, A(8) => 
                           out_b_8_port, A(7) => out_b_7_port, A(6) => 
                           out_b_6_port, A(5) => out_b_5_port, A(4) => 
                           out_b_4_port, A(3) => out_b_3_port, A(2) => 
                           out_b_2_port, A(1) => out_b_1_port, A(0) => 
                           out_b_0_port, B(31) => immediate_branch_31_port, 
                           B(30) => immediate_branch_30_port, B(29) => 
                           immediate_branch_29_port, B(28) => 
                           immediate_branch_28_port, B(27) => 
                           immediate_branch_27_port, B(26) => 
                           immediate_branch_26_port, B(25) => 
                           immediate_branch_25_port, B(24) => 
                           immediate_branch_24_port, B(23) => 
                           immediate_branch_23_port, B(22) => 
                           immediate_branch_22_port, B(21) => 
                           immediate_branch_21_port, B(20) => 
                           immediate_branch_20_port, B(19) => 
                           immediate_branch_19_port, B(18) => 
                           immediate_branch_18_port, B(17) => 
                           immediate_branch_17_port, B(16) => 
                           immediate_branch_16_port, B(15) => 
                           immediate_branch_15_port, B(14) => 
                           immediate_branch_14_port, B(13) => 
                           immediate_branch_13_port, B(12) => 
                           immediate_branch_12_port, B(11) => 
                           immediate_branch_11_port, B(10) => 
                           immediate_branch_10_port, B(9) => 
                           immediate_branch_9_port, B(8) => 
                           immediate_branch_8_port, B(7) => 
                           immediate_branch_7_port, B(6) => 
                           immediate_branch_6_port, B(5) => 
                           immediate_branch_5_port, B(4) => 
                           immediate_branch_4_port, B(3) => 
                           immediate_branch_3_port, B(2) => 
                           immediate_branch_2_port, B(1) => 
                           immediate_branch_1_port, B(0) => 
                           immediate_branch_0_port, SEL => S2, Y(31) => 
                           out_mux_2_31_port, Y(30) => out_mux_2_30_port, Y(29)
                           => out_mux_2_29_port, Y(28) => out_mux_2_28_port, 
                           Y(27) => out_mux_2_27_port, Y(26) => 
                           out_mux_2_26_port, Y(25) => out_mux_2_25_port, Y(24)
                           => out_mux_2_24_port, Y(23) => out_mux_2_23_port, 
                           Y(22) => out_mux_2_22_port, Y(21) => 
                           out_mux_2_21_port, Y(20) => out_mux_2_20_port, Y(19)
                           => out_mux_2_19_port, Y(18) => out_mux_2_18_port, 
                           Y(17) => out_mux_2_17_port, Y(16) => 
                           out_mux_2_16_port, Y(15) => out_mux_2_15_port, Y(14)
                           => out_mux_2_14_port, Y(13) => out_mux_2_13_port, 
                           Y(12) => out_mux_2_12_port, Y(11) => 
                           out_mux_2_11_port, Y(10) => out_mux_2_10_port, Y(9) 
                           => out_mux_2_9_port, Y(8) => out_mux_2_8_port, Y(7) 
                           => out_mux_2_7_port, Y(6) => out_mux_2_6_port, Y(5) 
                           => out_mux_2_5_port, Y(4) => out_mux_2_4_port, Y(3) 
                           => out_mux_2_3_port, Y(2) => out_mux_2_2_port, Y(1) 
                           => out_mux_2_1_port, Y(0) => out_mux_2_0_port);
   alu_dlx : ALU_N32 port map( AluOpCode(2) => aluopcode_i_2_port, AluOpCode(1)
                           => aluopcode_i_1_port, AluOpCode(0) => 
                           aluopcode_i_0_port, CompareOpCode(3) => 
                           compare_code_i_3_port, CompareOpCode(2) => 
                           compare_code_i_2_port, CompareOpCode(1) => 
                           compare_code_i_1_port, CompareOpCode(0) => 
                           compare_code_i_0_port, Add_subn => add_sub_i, 
                           ShiftOpCode(2) => shiftopcode_i_2_port, 
                           ShiftOpCode(1) => shiftopcode_i_1_port, 
                           ShiftOpCode(0) => shiftopcode_i_0_port, DATA1(31) =>
                           out_mux_1_31_port, DATA1(30) => out_mux_1_30_port, 
                           DATA1(29) => out_mux_1_29_port, DATA1(28) => 
                           out_mux_1_28_port, DATA1(27) => out_mux_1_27_port, 
                           DATA1(26) => out_mux_1_26_port, DATA1(25) => 
                           out_mux_1_25_port, DATA1(24) => out_mux_1_24_port, 
                           DATA1(23) => out_mux_1_23_port, DATA1(22) => 
                           out_mux_1_22_port, DATA1(21) => out_mux_1_21_port, 
                           DATA1(20) => out_mux_1_20_port, DATA1(19) => 
                           out_mux_1_19_port, DATA1(18) => out_mux_1_18_port, 
                           DATA1(17) => out_mux_1_17_port, DATA1(16) => 
                           out_mux_1_16_port, DATA1(15) => out_mux_1_15_port, 
                           DATA1(14) => out_mux_1_14_port, DATA1(13) => 
                           out_mux_1_13_port, DATA1(12) => out_mux_1_12_port, 
                           DATA1(11) => out_mux_1_11_port, DATA1(10) => 
                           out_mux_1_10_port, DATA1(9) => out_mux_1_9_port, 
                           DATA1(8) => out_mux_1_8_port, DATA1(7) => 
                           out_mux_1_7_port, DATA1(6) => out_mux_1_6_port, 
                           DATA1(5) => out_mux_1_5_port, DATA1(4) => 
                           out_mux_1_4_port, DATA1(3) => out_mux_1_3_port, 
                           DATA1(2) => out_mux_1_2_port, DATA1(1) => 
                           out_mux_1_1_port, DATA1(0) => out_mux_1_0_port, 
                           DATA2(31) => out_mux_2_31_port, DATA2(30) => 
                           out_mux_2_30_port, DATA2(29) => out_mux_2_29_port, 
                           DATA2(28) => out_mux_2_28_port, DATA2(27) => 
                           out_mux_2_27_port, DATA2(26) => out_mux_2_26_port, 
                           DATA2(25) => out_mux_2_25_port, DATA2(24) => 
                           out_mux_2_24_port, DATA2(23) => out_mux_2_23_port, 
                           DATA2(22) => out_mux_2_22_port, DATA2(21) => 
                           out_mux_2_21_port, DATA2(20) => out_mux_2_20_port, 
                           DATA2(19) => out_mux_2_19_port, DATA2(18) => 
                           out_mux_2_18_port, DATA2(17) => out_mux_2_17_port, 
                           DATA2(16) => out_mux_2_16_port, DATA2(15) => 
                           out_mux_2_15_port, DATA2(14) => out_mux_2_14_port, 
                           DATA2(13) => out_mux_2_13_port, DATA2(12) => 
                           out_mux_2_12_port, DATA2(11) => out_mux_2_11_port, 
                           DATA2(10) => out_mux_2_10_port, DATA2(9) => 
                           out_mux_2_9_port, DATA2(8) => out_mux_2_8_port, 
                           DATA2(7) => out_mux_2_7_port, DATA2(6) => 
                           out_mux_2_6_port, DATA2(5) => out_mux_2_5_port, 
                           DATA2(4) => out_mux_2_4_port, DATA2(3) => 
                           out_mux_2_3_port, DATA2(2) => out_mux_2_2_port, 
                           DATA2(1) => out_mux_2_1_port, DATA2(0) => 
                           out_mux_2_0_port, OUTALU(31) => reg_alu_in_31_port, 
                           OUTALU(30) => reg_alu_in_30_port, OUTALU(29) => 
                           reg_alu_in_29_port, OUTALU(28) => reg_alu_in_28_port
                           , OUTALU(27) => reg_alu_in_27_port, OUTALU(26) => 
                           reg_alu_in_26_port, OUTALU(25) => reg_alu_in_25_port
                           , OUTALU(24) => reg_alu_in_24_port, OUTALU(23) => 
                           reg_alu_in_23_port, OUTALU(22) => reg_alu_in_22_port
                           , OUTALU(21) => reg_alu_in_21_port, OUTALU(20) => 
                           reg_alu_in_20_port, OUTALU(19) => reg_alu_in_19_port
                           , OUTALU(18) => reg_alu_in_18_port, OUTALU(17) => 
                           reg_alu_in_17_port, OUTALU(16) => reg_alu_in_16_port
                           , OUTALU(15) => reg_alu_in_15_port, OUTALU(14) => 
                           reg_alu_in_14_port, OUTALU(13) => reg_alu_in_13_port
                           , OUTALU(12) => reg_alu_in_12_port, OUTALU(11) => 
                           reg_alu_in_11_port, OUTALU(10) => reg_alu_in_10_port
                           , OUTALU(9) => reg_alu_in_9_port, OUTALU(8) => 
                           reg_alu_in_8_port, OUTALU(7) => reg_alu_in_7_port, 
                           OUTALU(6) => reg_alu_in_6_port, OUTALU(5) => 
                           reg_alu_in_5_port, OUTALU(4) => reg_alu_in_4_port, 
                           OUTALU(3) => reg_alu_in_3_port, OUTALU(2) => 
                           reg_alu_in_2_port, OUTALU(1) => reg_alu_in_1_port, 
                           OUTALU(0) => reg_alu_in_0_port, return_address(31) 
                           => return_alu_31_port, return_address(30) => 
                           return_alu_30_port, return_address(29) => 
                           return_alu_29_port, return_address(28) => 
                           return_alu_28_port, return_address(27) => 
                           return_alu_27_port, return_address(26) => 
                           return_alu_26_port, return_address(25) => 
                           return_alu_25_port, return_address(24) => 
                           return_alu_24_port, return_address(23) => 
                           return_alu_23_port, return_address(22) => 
                           return_alu_22_port, return_address(21) => 
                           return_alu_21_port, return_address(20) => 
                           return_alu_20_port, return_address(19) => 
                           return_alu_19_port, return_address(18) => 
                           return_alu_18_port, return_address(17) => 
                           return_alu_17_port, return_address(16) => 
                           return_alu_16_port, return_address(15) => 
                           return_alu_15_port, return_address(14) => 
                           return_alu_14_port, return_address(13) => 
                           return_alu_13_port, return_address(12) => 
                           return_alu_12_port, return_address(11) => 
                           return_alu_11_port, return_address(10) => 
                           return_alu_10_port, return_address(9) => 
                           return_alu_9_port, return_address(8) => 
                           return_alu_8_port, return_address(7) => 
                           return_alu_7_port, return_address(6) => 
                           return_alu_6_port, return_address(5) => 
                           return_alu_5_port, return_address(4) => 
                           return_alu_4_port, return_address(3) => 
                           return_alu_3_port, return_address(2) => 
                           return_alu_2_port, return_address(1) => 
                           return_alu_1_port, return_address(0) => 
                           return_alu_0_port, CompBranch => comp_branch_i);
   alu_opcode_generator : AluOpCodeGen port map( IR_opcode(5) => 
                           aluopcode_reg_out_16_port, IR_opcode(4) => 
                           aluopcode_reg_out_15_port, IR_opcode(3) => 
                           aluopcode_reg_out_14_port, IR_opcode(2) => 
                           aluopcode_reg_out_13_port, IR_opcode(1) => 
                           aluopcode_reg_out_12_port, IR_opcode(0) => 
                           aluopcode_reg_out_11_port, IR_func(10) => 
                           aluopcode_reg_out_10_port, IR_func(9) => 
                           aluopcode_reg_out_9_port, IR_func(8) => 
                           aluopcode_reg_out_8_port, IR_func(7) => 
                           aluopcode_reg_out_7_port, IR_func(6) => 
                           aluopcode_reg_out_6_port, IR_func(5) => 
                           aluopcode_reg_out_5_port, IR_func(4) => 
                           aluopcode_reg_out_4_port, IR_func(3) => 
                           aluopcode_reg_out_3_port, IR_func(2) => 
                           aluopcode_reg_out_2_port, IR_func(1) => 
                           aluopcode_reg_out_1_port, IR_func(0) => 
                           aluopcode_reg_out_0_port, AluOpCode(2) => 
                           aluopcode_i_2_port, AluOpCode(1) => 
                           aluopcode_i_1_port, AluOpCode(0) => 
                           aluopcode_i_0_port, Add_Subn => add_sub_i, 
                           CompareCode(3) => compare_code_i_3_port, 
                           CompareCode(2) => compare_code_i_2_port, 
                           CompareCode(1) => compare_code_i_1_port, 
                           CompareCode(0) => compare_code_i_0_port, 
                           ShiftOpCode(2) => shiftopcode_i_2_port, 
                           ShiftOpCode(1) => shiftopcode_i_1_port, 
                           ShiftOpCode(0) => shiftopcode_i_0_port);
   reg_alu_out : registro_N32_5 port map( data(31) => reg_alu_in_31_port, 
                           data(30) => reg_alu_in_30_port, data(29) => 
                           reg_alu_in_29_port, data(28) => reg_alu_in_28_port, 
                           data(27) => reg_alu_in_27_port, data(26) => 
                           reg_alu_in_26_port, data(25) => reg_alu_in_25_port, 
                           data(24) => reg_alu_in_24_port, data(23) => 
                           reg_alu_in_23_port, data(22) => reg_alu_in_22_port, 
                           data(21) => reg_alu_in_21_port, data(20) => 
                           reg_alu_in_20_port, data(19) => reg_alu_in_19_port, 
                           data(18) => reg_alu_in_18_port, data(17) => 
                           reg_alu_in_17_port, data(16) => reg_alu_in_16_port, 
                           data(15) => reg_alu_in_15_port, data(14) => 
                           reg_alu_in_14_port, data(13) => reg_alu_in_13_port, 
                           data(12) => reg_alu_in_12_port, data(11) => 
                           reg_alu_in_11_port, data(10) => reg_alu_in_10_port, 
                           data(9) => reg_alu_in_9_port, data(8) => 
                           reg_alu_in_8_port, data(7) => reg_alu_in_7_port, 
                           data(6) => reg_alu_in_6_port, data(5) => 
                           reg_alu_in_5_port, data(4) => reg_alu_in_4_port, 
                           data(3) => reg_alu_in_3_port, data(2) => 
                           reg_alu_in_2_port, data(1) => reg_alu_in_1_port, 
                           data(0) => reg_alu_in_0_port, enable => EN_regOUTALU
                           , clock => clk, clear => rst, Q(31) => 
                           ADD_mem_31_port, Q(30) => ADD_mem_30_port, Q(29) => 
                           ADD_mem_29_port, Q(28) => ADD_mem_28_port, Q(27) => 
                           ADD_mem_27_port, Q(26) => ADD_mem_26_port, Q(25) => 
                           ADD_mem_25_port, Q(24) => ADD_mem_24_port, Q(23) => 
                           ADD_mem_23_port, Q(22) => ADD_mem_22_port, Q(21) => 
                           ADD_mem_21_port, Q(20) => ADD_mem_20_port, Q(19) => 
                           ADD_mem_19_port, Q(18) => ADD_mem_18_port, Q(17) => 
                           ADD_mem_17_port, Q(16) => ADD_mem_16_port, Q(15) => 
                           ADD_mem_15_port, Q(14) => ADD_mem_14_port, Q(13) => 
                           ADD_mem_13_port, Q(12) => ADD_mem_12_port, Q(11) => 
                           ADD_mem_11_port, Q(10) => ADD_mem_10_port, Q(9) => 
                           ADD_mem_9_port, Q(8) => ADD_mem_8_port, Q(7) => 
                           ADD_mem_7_port, Q(6) => ADD_mem_6_port, Q(5) => 
                           ADD_mem_5_port, Q(4) => ADD_mem_4_port, Q(3) => 
                           ADD_mem_3_port, Q(2) => ADD_mem_2_port, Q(1) => 
                           ADD_mem_1_port, Q(0) => ADD_mem_0_port);
   reg_b2 : registro_N32_4 port map( data(31) => out_b_31_port, data(30) => 
                           out_b_30_port, data(29) => out_b_29_port, data(28) 
                           => out_b_28_port, data(27) => out_b_27_port, 
                           data(26) => out_b_26_port, data(25) => out_b_25_port
                           , data(24) => out_b_24_port, data(23) => 
                           out_b_23_port, data(22) => out_b_22_port, data(21) 
                           => out_b_21_port, data(20) => out_b_20_port, 
                           data(19) => out_b_19_port, data(18) => out_b_18_port
                           , data(17) => out_b_17_port, data(16) => 
                           out_b_16_port, data(15) => out_b_15_port, data(14) 
                           => out_b_14_port, data(13) => out_b_13_port, 
                           data(12) => out_b_12_port, data(11) => out_b_11_port
                           , data(10) => out_b_10_port, data(9) => out_b_9_port
                           , data(8) => out_b_8_port, data(7) => out_b_7_port, 
                           data(6) => out_b_6_port, data(5) => out_b_5_port, 
                           data(4) => out_b_4_port, data(3) => out_b_3_port, 
                           data(2) => out_b_2_port, data(1) => out_b_1_port, 
                           data(0) => out_b_0_port, enable => EN_regB2, clock 
                           => clk, clear => rst, Q(31) => DIN_mem(31), Q(30) =>
                           DIN_mem(30), Q(29) => DIN_mem(29), Q(28) => 
                           DIN_mem(28), Q(27) => DIN_mem(27), Q(26) => 
                           DIN_mem(26), Q(25) => DIN_mem(25), Q(24) => 
                           DIN_mem(24), Q(23) => DIN_mem(23), Q(22) => 
                           DIN_mem(22), Q(21) => DIN_mem(21), Q(20) => 
                           DIN_mem(20), Q(19) => DIN_mem(19), Q(18) => 
                           DIN_mem(18), Q(17) => DIN_mem(17), Q(16) => 
                           DIN_mem(16), Q(15) => DIN_mem(15), Q(14) => 
                           DIN_mem(14), Q(13) => DIN_mem(13), Q(12) => 
                           DIN_mem(12), Q(11) => DIN_mem(11), Q(10) => 
                           DIN_mem(10), Q(9) => DIN_mem(9), Q(8) => DIN_mem(8),
                           Q(7) => DIN_mem(7), Q(6) => DIN_mem(6), Q(5) => 
                           DIN_mem(5), Q(4) => DIN_mem(4), Q(3) => DIN_mem(3), 
                           Q(2) => DIN_mem(2), Q(1) => DIN_mem(1), Q(0) => 
                           DIN_mem(0));
   reg_rd2 : registro_N5_2 port map( data(4) => out_rd1_4_port, data(3) => 
                           out_rd1_3_port, data(2) => out_rd1_2_port, data(1) 
                           => out_rd1_1_port, data(0) => out_rd1_0_port, enable
                           => EN_regRD2, clock => clk, clear => rst, Q(4) => 
                           out_rd2_4_port, Q(3) => out_rd2_3_port, Q(2) => 
                           out_rd2_2_port, Q(1) => out_rd2_1_port, Q(0) => 
                           out_rd2_0_port);
   reg_return : registro_N32_3 port map( data(31) => return_alu_31_port, 
                           data(30) => return_alu_30_port, data(29) => 
                           return_alu_29_port, data(28) => return_alu_28_port, 
                           data(27) => return_alu_27_port, data(26) => 
                           return_alu_26_port, data(25) => return_alu_25_port, 
                           data(24) => return_alu_24_port, data(23) => 
                           return_alu_23_port, data(22) => return_alu_22_port, 
                           data(21) => return_alu_21_port, data(20) => 
                           return_alu_20_port, data(19) => return_alu_19_port, 
                           data(18) => return_alu_18_port, data(17) => 
                           return_alu_17_port, data(16) => return_alu_16_port, 
                           data(15) => return_alu_15_port, data(14) => 
                           return_alu_14_port, data(13) => return_alu_13_port, 
                           data(12) => return_alu_12_port, data(11) => 
                           return_alu_11_port, data(10) => return_alu_10_port, 
                           data(9) => return_alu_9_port, data(8) => 
                           return_alu_8_port, data(7) => return_alu_7_port, 
                           data(6) => return_alu_6_port, data(5) => 
                           return_alu_5_port, data(4) => return_alu_4_port, 
                           data(3) => return_alu_3_port, data(2) => 
                           return_alu_2_port, data(1) => return_alu_1_port, 
                           data(0) => return_alu_0_port, enable => EN_regRET, 
                           clock => clk, clear => rst, Q(31) => 
                           return_out_31_port, Q(30) => return_out_30_port, 
                           Q(29) => return_out_29_port, Q(28) => 
                           return_out_28_port, Q(27) => return_out_27_port, 
                           Q(26) => return_out_26_port, Q(25) => 
                           return_out_25_port, Q(24) => return_out_24_port, 
                           Q(23) => return_out_23_port, Q(22) => 
                           return_out_22_port, Q(21) => return_out_21_port, 
                           Q(20) => return_out_20_port, Q(19) => 
                           return_out_19_port, Q(18) => return_out_18_port, 
                           Q(17) => return_out_17_port, Q(16) => 
                           return_out_16_port, Q(15) => return_out_15_port, 
                           Q(14) => return_out_14_port, Q(13) => 
                           return_out_13_port, Q(12) => return_out_12_port, 
                           Q(11) => return_out_11_port, Q(10) => 
                           return_out_10_port, Q(9) => return_out_9_port, Q(8) 
                           => return_out_8_port, Q(7) => return_out_7_port, 
                           Q(6) => return_out_6_port, Q(5) => return_out_5_port
                           , Q(4) => return_out_4_port, Q(3) => 
                           return_out_3_port, Q(2) => return_out_2_port, Q(1) 
                           => return_out_1_port, Q(0) => return_out_0_port);
   mux_ret_alu : mux21_N32_2 port map( A(31) => ADD_mem_31_port, A(30) => 
                           ADD_mem_30_port, A(29) => ADD_mem_29_port, A(28) => 
                           ADD_mem_28_port, A(27) => ADD_mem_27_port, A(26) => 
                           ADD_mem_26_port, A(25) => ADD_mem_25_port, A(24) => 
                           ADD_mem_24_port, A(23) => ADD_mem_23_port, A(22) => 
                           ADD_mem_22_port, A(21) => ADD_mem_21_port, A(20) => 
                           ADD_mem_20_port, A(19) => ADD_mem_19_port, A(18) => 
                           ADD_mem_18_port, A(17) => ADD_mem_17_port, A(16) => 
                           ADD_mem_16_port, A(15) => ADD_mem_15_port, A(14) => 
                           ADD_mem_14_port, A(13) => ADD_mem_13_port, A(12) => 
                           ADD_mem_12_port, A(11) => ADD_mem_11_port, A(10) => 
                           ADD_mem_10_port, A(9) => ADD_mem_9_port, A(8) => 
                           ADD_mem_8_port, A(7) => ADD_mem_7_port, A(6) => 
                           ADD_mem_6_port, A(5) => ADD_mem_5_port, A(4) => 
                           ADD_mem_4_port, A(3) => ADD_mem_3_port, A(2) => 
                           ADD_mem_2_port, A(1) => ADD_mem_1_port, A(0) => 
                           ADD_mem_0_port, B(31) => return_out_31_port, B(30) 
                           => return_out_30_port, B(29) => return_out_29_port, 
                           B(28) => return_out_28_port, B(27) => 
                           return_out_27_port, B(26) => return_out_26_port, 
                           B(25) => return_out_25_port, B(24) => 
                           return_out_24_port, B(23) => return_out_23_port, 
                           B(22) => return_out_22_port, B(21) => 
                           return_out_21_port, B(20) => return_out_20_port, 
                           B(19) => return_out_19_port, B(18) => 
                           return_out_18_port, B(17) => return_out_17_port, 
                           B(16) => return_out_16_port, B(15) => 
                           return_out_15_port, B(14) => return_out_14_port, 
                           B(13) => return_out_13_port, B(12) => 
                           return_out_12_port, B(11) => return_out_11_port, 
                           B(10) => return_out_10_port, B(9) => 
                           return_out_9_port, B(8) => return_out_8_port, B(7) 
                           => return_out_7_port, B(6) => return_out_6_port, 
                           B(5) => return_out_5_port, B(4) => return_out_4_port
                           , B(3) => return_out_3_port, B(2) => 
                           return_out_2_port, B(1) => return_out_1_port, B(0) 
                           => return_out_0_port, SEL => Sel_ret_alu, Y(31) => 
                           out_ret_alu_31_port, Y(30) => out_ret_alu_30_port, 
                           Y(29) => out_ret_alu_29_port, Y(28) => 
                           out_ret_alu_28_port, Y(27) => out_ret_alu_27_port, 
                           Y(26) => out_ret_alu_26_port, Y(25) => 
                           out_ret_alu_25_port, Y(24) => out_ret_alu_24_port, 
                           Y(23) => out_ret_alu_23_port, Y(22) => 
                           out_ret_alu_22_port, Y(21) => out_ret_alu_21_port, 
                           Y(20) => out_ret_alu_20_port, Y(19) => 
                           out_ret_alu_19_port, Y(18) => out_ret_alu_18_port, 
                           Y(17) => out_ret_alu_17_port, Y(16) => 
                           out_ret_alu_16_port, Y(15) => out_ret_alu_15_port, 
                           Y(14) => out_ret_alu_14_port, Y(13) => 
                           out_ret_alu_13_port, Y(12) => out_ret_alu_12_port, 
                           Y(11) => out_ret_alu_11_port, Y(10) => 
                           out_ret_alu_10_port, Y(9) => out_ret_alu_9_port, 
                           Y(8) => out_ret_alu_8_port, Y(7) => 
                           out_ret_alu_7_port, Y(6) => out_ret_alu_6_port, Y(5)
                           => out_ret_alu_5_port, Y(4) => out_ret_alu_4_port, 
                           Y(3) => out_ret_alu_3_port, Y(2) => 
                           out_ret_alu_2_port, Y(1) => out_ret_alu_1_port, Y(0)
                           => out_ret_alu_0_port);
   reg_alu2 : registro_N32_2 port map( data(31) => out_ret_alu_31_port, 
                           data(30) => out_ret_alu_30_port, data(29) => 
                           out_ret_alu_29_port, data(28) => out_ret_alu_28_port
                           , data(27) => out_ret_alu_27_port, data(26) => 
                           out_ret_alu_26_port, data(25) => out_ret_alu_25_port
                           , data(24) => out_ret_alu_24_port, data(23) => 
                           out_ret_alu_23_port, data(22) => out_ret_alu_22_port
                           , data(21) => out_ret_alu_21_port, data(20) => 
                           out_ret_alu_20_port, data(19) => out_ret_alu_19_port
                           , data(18) => out_ret_alu_18_port, data(17) => 
                           out_ret_alu_17_port, data(16) => out_ret_alu_16_port
                           , data(15) => out_ret_alu_15_port, data(14) => 
                           out_ret_alu_14_port, data(13) => out_ret_alu_13_port
                           , data(12) => out_ret_alu_12_port, data(11) => 
                           out_ret_alu_11_port, data(10) => out_ret_alu_10_port
                           , data(9) => out_ret_alu_9_port, data(8) => 
                           out_ret_alu_8_port, data(7) => out_ret_alu_7_port, 
                           data(6) => out_ret_alu_6_port, data(5) => 
                           out_ret_alu_5_port, data(4) => out_ret_alu_4_port, 
                           data(3) => out_ret_alu_3_port, data(2) => 
                           out_ret_alu_2_port, data(1) => out_ret_alu_1_port, 
                           data(0) => out_ret_alu_0_port, enable => EN_regALU2,
                           clock => clk, clear => rst, Q(31) => alu2_31_port, 
                           Q(30) => alu2_30_port, Q(29) => alu2_29_port, Q(28) 
                           => alu2_28_port, Q(27) => alu2_27_port, Q(26) => 
                           alu2_26_port, Q(25) => alu2_25_port, Q(24) => 
                           alu2_24_port, Q(23) => alu2_23_port, Q(22) => 
                           alu2_22_port, Q(21) => alu2_21_port, Q(20) => 
                           alu2_20_port, Q(19) => alu2_19_port, Q(18) => 
                           alu2_18_port, Q(17) => alu2_17_port, Q(16) => 
                           alu2_16_port, Q(15) => alu2_15_port, Q(14) => 
                           alu2_14_port, Q(13) => alu2_13_port, Q(12) => 
                           alu2_12_port, Q(11) => alu2_11_port, Q(10) => 
                           alu2_10_port, Q(9) => alu2_9_port, Q(8) => 
                           alu2_8_port, Q(7) => alu2_7_port, Q(6) => 
                           alu2_6_port, Q(5) => alu2_5_port, Q(4) => 
                           alu2_4_port, Q(3) => alu2_3_port, Q(2) => 
                           alu2_2_port, Q(1) => alu2_1_port, Q(0) => 
                           alu2_0_port);
   reg_lmd : registro_N32_1 port map( data(31) => DOUT_mem(31), data(30) => 
                           DOUT_mem(30), data(29) => DOUT_mem(29), data(28) => 
                           DOUT_mem(28), data(27) => DOUT_mem(27), data(26) => 
                           DOUT_mem(26), data(25) => DOUT_mem(25), data(24) => 
                           DOUT_mem(24), data(23) => DOUT_mem(23), data(22) => 
                           DOUT_mem(22), data(21) => DOUT_mem(21), data(20) => 
                           DOUT_mem(20), data(19) => DOUT_mem(19), data(18) => 
                           DOUT_mem(18), data(17) => DOUT_mem(17), data(16) => 
                           DOUT_mem(16), data(15) => DOUT_mem(15), data(14) => 
                           DOUT_mem(14), data(13) => DOUT_mem(13), data(12) => 
                           DOUT_mem(12), data(11) => DOUT_mem(11), data(10) => 
                           DOUT_mem(10), data(9) => DOUT_mem(9), data(8) => 
                           DOUT_mem(8), data(7) => DOUT_mem(7), data(6) => 
                           DOUT_mem(6), data(5) => DOUT_mem(5), data(4) => 
                           DOUT_mem(4), data(3) => DOUT_mem(3), data(2) => 
                           DOUT_mem(2), data(1) => DOUT_mem(1), data(0) => 
                           DOUT_mem(0), enable => EN_regLMD, clock => clk, 
                           clear => rst, Q(31) => lmd_31_port, Q(30) => 
                           lmd_30_port, Q(29) => lmd_29_port, Q(28) => 
                           lmd_28_port, Q(27) => lmd_27_port, Q(26) => 
                           lmd_26_port, Q(25) => lmd_25_port, Q(24) => 
                           lmd_24_port, Q(23) => lmd_23_port, Q(22) => 
                           lmd_22_port, Q(21) => lmd_21_port, Q(20) => 
                           lmd_20_port, Q(19) => lmd_19_port, Q(18) => 
                           lmd_18_port, Q(17) => lmd_17_port, Q(16) => 
                           lmd_16_port, Q(15) => lmd_15_port, Q(14) => 
                           lmd_14_port, Q(13) => lmd_13_port, Q(12) => 
                           lmd_12_port, Q(11) => lmd_11_port, Q(10) => 
                           lmd_10_port, Q(9) => lmd_9_port, Q(8) => lmd_8_port,
                           Q(7) => lmd_7_port, Q(6) => lmd_6_port, Q(5) => 
                           lmd_5_port, Q(4) => lmd_4_port, Q(3) => lmd_3_port, 
                           Q(2) => lmd_2_port, Q(1) => lmd_1_port, Q(0) => 
                           lmd_0_port);
   reg_rd3 : registro_N5_1 port map( data(4) => out_rd2_4_port, data(3) => 
                           out_rd2_3_port, data(2) => out_rd2_2_port, data(1) 
                           => out_rd2_1_port, data(0) => out_rd2_0_port, enable
                           => EN_regRD3, clock => clk, clear => rst, Q(4) => 
                           rd3_4_port, Q(3) => rd3_3_port, Q(2) => rd3_2_port, 
                           Q(1) => rd3_1_port, Q(0) => rd3_0_port);
   mux_lmd_alu : mux21_N32_1 port map( A(31) => alu2_31_port, A(30) => 
                           alu2_30_port, A(29) => alu2_29_port, A(28) => 
                           alu2_28_port, A(27) => alu2_27_port, A(26) => 
                           alu2_26_port, A(25) => alu2_25_port, A(24) => 
                           alu2_24_port, A(23) => alu2_23_port, A(22) => 
                           alu2_22_port, A(21) => alu2_21_port, A(20) => 
                           alu2_20_port, A(19) => alu2_19_port, A(18) => 
                           alu2_18_port, A(17) => alu2_17_port, A(16) => 
                           alu2_16_port, A(15) => alu2_15_port, A(14) => 
                           alu2_14_port, A(13) => alu2_13_port, A(12) => 
                           alu2_12_port, A(11) => alu2_11_port, A(10) => 
                           alu2_10_port, A(9) => alu2_9_port, A(8) => 
                           alu2_8_port, A(7) => alu2_7_port, A(6) => 
                           alu2_6_port, A(5) => alu2_5_port, A(4) => 
                           alu2_4_port, A(3) => alu2_3_port, A(2) => 
                           alu2_2_port, A(1) => alu2_1_port, A(0) => 
                           alu2_0_port, B(31) => lmd_31_port, B(30) => 
                           lmd_30_port, B(29) => lmd_29_port, B(28) => 
                           lmd_28_port, B(27) => lmd_27_port, B(26) => 
                           lmd_26_port, B(25) => lmd_25_port, B(24) => 
                           lmd_24_port, B(23) => lmd_23_port, B(22) => 
                           lmd_22_port, B(21) => lmd_21_port, B(20) => 
                           lmd_20_port, B(19) => lmd_19_port, B(18) => 
                           lmd_18_port, B(17) => lmd_17_port, B(16) => 
                           lmd_16_port, B(15) => lmd_15_port, B(14) => 
                           lmd_14_port, B(13) => lmd_13_port, B(12) => 
                           lmd_12_port, B(11) => lmd_11_port, B(10) => 
                           lmd_10_port, B(9) => lmd_9_port, B(8) => lmd_8_port,
                           B(7) => lmd_7_port, B(6) => lmd_6_port, B(5) => 
                           lmd_5_port, B(4) => lmd_4_port, B(3) => lmd_3_port, 
                           B(2) => lmd_2_port, B(1) => lmd_1_port, B(0) => 
                           lmd_0_port, SEL => Sel_alu_lmd, Y(31) => 
                           alu2_lmd_31_port, Y(30) => alu2_lmd_30_port, Y(29) 
                           => alu2_lmd_29_port, Y(28) => alu2_lmd_28_port, 
                           Y(27) => alu2_lmd_27_port, Y(26) => alu2_lmd_26_port
                           , Y(25) => alu2_lmd_25_port, Y(24) => 
                           alu2_lmd_24_port, Y(23) => alu2_lmd_23_port, Y(22) 
                           => alu2_lmd_22_port, Y(21) => alu2_lmd_21_port, 
                           Y(20) => alu2_lmd_20_port, Y(19) => alu2_lmd_19_port
                           , Y(18) => alu2_lmd_18_port, Y(17) => 
                           alu2_lmd_17_port, Y(16) => alu2_lmd_16_port, Y(15) 
                           => alu2_lmd_15_port, Y(14) => alu2_lmd_14_port, 
                           Y(13) => alu2_lmd_13_port, Y(12) => alu2_lmd_12_port
                           , Y(11) => alu2_lmd_11_port, Y(10) => 
                           alu2_lmd_10_port, Y(9) => alu2_lmd_9_port, Y(8) => 
                           alu2_lmd_8_port, Y(7) => alu2_lmd_7_port, Y(6) => 
                           alu2_lmd_6_port, Y(5) => alu2_lmd_5_port, Y(4) => 
                           alu2_lmd_4_port, Y(3) => alu2_lmd_3_port, Y(2) => 
                           alu2_lmd_2_port, Y(1) => alu2_lmd_1_port, Y(0) => 
                           alu2_lmd_0_port);
   mux_address_write : mux21_N5 port map( A(4) => rd3_4_port, A(3) => 
                           rd3_3_port, A(2) => rd3_2_port, A(1) => rd3_1_port, 
                           A(0) => rd3_0_port, B(4) => X_Logic1_port, B(3) => 
                           X_Logic1_port, B(2) => X_Logic1_port, B(1) => 
                           X_Logic1_port, B(0) => X_Logic1_port, SEL => 
                           sel_31_rd, Y(4) => add_w_rf_4_port, Y(3) => 
                           add_w_rf_3_port, Y(2) => add_w_rf_2_port, Y(1) => 
                           add_w_rf_1_port, Y(0) => add_w_rf_0_port);
   U3 : CLKBUF_X3 port map( A => reset_pipe2, Z => n1);
   U4 : NOR4_X2 port map( A1 => IR_dp(26), A2 => n8, A3 => IR_dp(28), A4 => 
                           IR_dp(27), ZN => n7);
   U5 : NOR2_X1 port map( A1 => flush, A2 => n2, ZN => reset_pipe2);
   U6 : INV_X1 port map( A => rst, ZN => n2);
   U7 : NAND2_X1 port map( A1 => n3, A2 => n4, ZN => N56);
   U8 : NAND3_X1 port map( A1 => n5, A2 => n6, A3 => IR_dp(28), ZN => n4);
   U9 : INV_X1 port map( A => N40, ZN => n3);
   U10 : MUX2_X1 port map( A => IR_dp(20), B => IR_dp(15), S => n7, Z => N55);
   U11 : MUX2_X1 port map( A => IR_dp(19), B => IR_dp(14), S => n7, Z => N53);
   U12 : MUX2_X1 port map( A => IR_dp(18), B => IR_dp(13), S => n7, Z => N51);
   U13 : MUX2_X1 port map( A => IR_dp(17), B => IR_dp(12), S => n7, Z => N49);
   U14 : MUX2_X1 port map( A => IR_dp(16), B => IR_dp(11), S => n7, Z => N47);
   U15 : NOR3_X1 port map( A1 => n8, A2 => IR_dp(28), A3 => n6, ZN => N40);
   U16 : INV_X1 port map( A => IR_dp(27), ZN => n6);
   U17 : INV_X1 port map( A => n5, ZN => n8);
   U18 : NOR3_X1 port map( A1 => IR_dp(31), A2 => IR_dp(30), A3 => IR_dp(29), 
                           ZN => n5);

end SYN_behaviour;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_DLX_IR_SIZE32_PC_SIZE32.all;

entity DLX_IR_SIZE32_PC_SIZE32 is

   port( Clk, Rst : in std_logic;  dram_RD, dram_WR : out std_logic;  dram_ADD,
         dram_DIN : out std_logic_vector (31 downto 0);  dram_DOUT : in 
         std_logic_vector (31 downto 0);  iram_Addr : out std_logic_vector (31 
         downto 0);  iram_Dout : in std_logic_vector (31 downto 0));

end DLX_IR_SIZE32_PC_SIZE32;

architecture SYN_dlx_rtl of DLX_IR_SIZE32_PC_SIZE32 is

   component NOR2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X2
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component AND2_X2
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component DLX_IR_SIZE32_PC_SIZE32_DW01_add_1
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component DLX_IR_SIZE32_PC_SIZE32_DW01_add_0
      port( A, B : in std_logic_vector (31 downto 0);  CI : in std_logic;  SUM 
            : out std_logic_vector (31 downto 0);  CO : out std_logic);
   end component;
   
   component 
      CU_HDW_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE21
      port( Clk, Rst : in std_logic;  IR_IN : in std_logic_vector (31 downto 0)
            ;  flush : in std_logic;  IR_LATCH_EN, NPC1_LATCH_EN, NPC2_LATCH_EN
            , RegA_LATCH_EN, RegB_LATCH_EN, RegAluOpCodeGen_EN, RegIMM_LATCH_EN
            , Reg_RD1_EN, RD1, RD2, B2_LATCH_EN, MUXA_SEL, MUXB_SEL, 
            ALU_OUTREG_EN, RETURN_REG_EN, Reg_RD2_EN, DRAM_WE, ALU_OUT2_SEL, 
            LMD_LATCH_EN, Alu_outreg2_en, JUMP_en, PC_LATCH_EN, Reg_RD3_EN, 
            write_stop_if_branch, WB_MUX_SEL, RF_WE, WB_MUX_ADD_SEL, WR : out 
            std_logic);
   end component;
   
   component mux21_N32_0
      port( A, B : in std_logic_vector (31 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (31 downto 0));
   end component;
   
   component datapath_reg_size32
      port( clk, rst, flush, RF1, RF2, WF1, EN_regA, EN_regB, EN_regIMM, 
            EN_regALUOP, EN_regRD1, EN_regNPC2, S1, S2, EN_regRET, EN_regOUTALU
            , EN_regB2, EN_regRD2, EN_regALU2, EN_regLMD, EN_regRD3, 
            Sel_ret_alu, Sel_alu_lmd, sel_31_rd : in std_logic;  NPC, IR_dp : 
            in std_logic_vector (31 downto 0);  OUT_DP : out std_logic_vector 
            (31 downto 0);  comp_branch_i : out std_logic;  immediate_branch, 
            ADD_mem, DIN_mem : out std_logic_vector (31 downto 0);  DOUT_mem : 
            in std_logic_vector (31 downto 0));
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal X_Logic1_port, X_Logic0_port, jump_verified, rd1_i, rd2_i, wr_i, 
      RegA_LATCH_EN_i, RegB_LATCH_EN_i, RegIMM_LATCH_EN_i, RegAluOpCodeGen_EN_i
      , en_RD1_i, NPC2_LATCH_EN_i, MUXA_SEL_i, MUXB_SEL_i, RETURN_REG_EN_i, 
      ALU_OUTREG_EN_i, B2_EN_i, en_RD2_i, Alu_outreg2_en_i, LMD_LATCH_EN_i, 
      en_RD3_i, sel_alu_ret_i, WB_MUX_SEL_i, wb_mux_add_sel_i, out_NPC_31_port,
      out_NPC_30_port, out_NPC_29_port, out_NPC_28_port, out_NPC_27_port, 
      out_NPC_26_port, out_NPC_25_port, out_NPC_24_port, out_NPC_23_port, 
      out_NPC_22_port, out_NPC_21_port, out_NPC_20_port, out_NPC_19_port, 
      out_NPC_18_port, out_NPC_17_port, out_NPC_16_port, out_NPC_15_port, 
      out_NPC_14_port, out_NPC_13_port, out_NPC_12_port, out_NPC_11_port, 
      out_NPC_10_port, out_NPC_9_port, out_NPC_8_port, out_NPC_7_port, 
      out_NPC_6_port, out_NPC_5_port, out_NPC_4_port, out_NPC_3_port, 
      out_NPC_2_port, out_NPC_1_port, out_NPC_0_port, IR_31_port, IR_30_port, 
      IR_29_port, IR_28_port, IR_27_port, IR_26_port, IR_25_port, IR_24_port, 
      IR_23_port, IR_22_port, IR_21_port, IR_20_port, IR_19_port, IR_18_port, 
      IR_17_port, IR_16_port, IR_15_port, IR_14_port, IR_13_port, IR_12_port, 
      IR_11_port, IR_10_port, IR_9_port, IR_8_port, IR_7_port, IR_6_port, 
      IR_5_port, IR_4_port, IR_3_port, IR_2_port, IR_1_port, IR_0_port, 
      comp_branch_dp, immediate_31_port, immediate_30_port, immediate_29_port, 
      immediate_28_port, immediate_27_port, immediate_26_port, 
      immediate_25_port, immediate_24_port, immediate_23_port, 
      immediate_22_port, immediate_21_port, immediate_20_port, 
      immediate_19_port, immediate_18_port, immediate_17_port, 
      immediate_16_port, immediate_15_port, immediate_14_port, 
      immediate_13_port, immediate_12_port, immediate_11_port, 
      immediate_10_port, immediate_9_port, immediate_8_port, immediate_7_port, 
      immediate_6_port, immediate_5_port, immediate_4_port, immediate_3_port, 
      immediate_2_port, immediate_1_port, immediate_0_port, PC_31_port, 
      PC_30_port, PC_29_port, PC_28_port, PC_27_port, PC_26_port, PC_25_port, 
      PC_24_port, PC_23_port, PC_22_port, PC_21_port, PC_20_port, PC_19_port, 
      PC_18_port, PC_17_port, PC_16_port, PC_15_port, PC_14_port, PC_13_port, 
      PC_12_port, PC_11_port, PC_10_port, PC_9_port, PC_8_port, PC_7_port, 
      PC_6_port, PC_5_port, PC_4_port, PC_3_port, PC_2_port, PC_1_port, 
      PC_0_port, PC_BUS_31_port, PC_BUS_30_port, PC_BUS_29_port, PC_BUS_28_port
      , PC_BUS_27_port, PC_BUS_26_port, PC_BUS_25_port, PC_BUS_24_port, 
      PC_BUS_23_port, PC_BUS_22_port, PC_BUS_21_port, PC_BUS_20_port, 
      PC_BUS_19_port, PC_BUS_18_port, PC_BUS_17_port, PC_BUS_16_port, 
      PC_BUS_15_port, PC_BUS_14_port, PC_BUS_13_port, PC_BUS_12_port, 
      PC_BUS_11_port, PC_BUS_10_port, PC_BUS_9_port, PC_BUS_8_port, 
      PC_BUS_7_port, PC_BUS_6_port, PC_BUS_5_port, PC_BUS_4_port, PC_BUS_3_port
      , PC_BUS_2_port, PC_BUS_1_port, PC_BUS_0_port, in_NPC_31_port, 
      in_NPC_30_port, in_NPC_29_port, in_NPC_28_port, in_NPC_27_port, 
      in_NPC_26_port, in_NPC_25_port, in_NPC_24_port, in_NPC_23_port, 
      in_NPC_22_port, in_NPC_21_port, in_NPC_20_port, in_NPC_19_port, 
      in_NPC_18_port, in_NPC_17_port, in_NPC_16_port, in_NPC_15_port, 
      in_NPC_14_port, in_NPC_13_port, in_NPC_12_port, in_NPC_11_port, 
      in_NPC_10_port, in_NPC_9_port, in_NPC_8_port, in_NPC_7_port, 
      in_NPC_6_port, in_NPC_5_port, in_NPC_4_port, in_NPC_3_port, in_NPC_2_port
      , in_NPC_1_port, in_NPC_0_port, NPC1_LATCH_EN_i, JUMP_EN_i, npc2_31_port,
      npc2_30_port, npc2_29_port, npc2_28_port, npc2_27_port, npc2_26_port, 
      npc2_25_port, npc2_24_port, npc2_23_port, npc2_22_port, npc2_21_port, 
      npc2_20_port, npc2_19_port, npc2_18_port, npc2_17_port, npc2_16_port, 
      npc2_15_port, npc2_14_port, npc2_13_port, npc2_12_port, npc2_11_port, 
      npc2_10_port, npc2_9_port, npc2_8_port, npc2_7_port, npc2_6_port, 
      npc2_5_port, npc2_4_port, npc2_3_port, npc2_2_port, npc2_1_port, 
      npc2_0_port, pc_jump_31_port, pc_jump_30_port, pc_jump_29_port, 
      pc_jump_28_port, pc_jump_27_port, pc_jump_26_port, pc_jump_25_port, 
      pc_jump_24_port, pc_jump_23_port, pc_jump_22_port, pc_jump_21_port, 
      pc_jump_20_port, pc_jump_19_port, pc_jump_18_port, pc_jump_17_port, 
      pc_jump_16_port, pc_jump_15_port, pc_jump_14_port, pc_jump_13_port, 
      pc_jump_12_port, pc_jump_11_port, pc_jump_10_port, pc_jump_9_port, 
      pc_jump_8_port, pc_jump_7_port, pc_jump_6_port, pc_jump_5_port, 
      pc_jump_4_port, pc_jump_3_port, pc_jump_2_port, pc_jump_1_port, 
      pc_jump_0_port, wr_cu, write_stop_if_branch_i, net583, net584, net585, 
      net714, net715, net716, net717, net718, net719, net720, net721, net722, 
      net723, net724, net725, net726, net727, net728, net729, net730, net731, 
      net732, net733, net734, net735, net736, net737, net738, net739, net740, 
      net741, net742, net743, net744, net745, n1, n2, net713, net712, net711, 
      net710, net709, net708, net707, net706, net705, net704, net703, net702, 
      net701, net700, net699, net698, net697, net696, net695, net694, net693, 
      net692, net691, net690, net689, net688, net687, net686, net685, net684, 
      net683, net682, net681, net680, net679, net678, net677, net676, net675, 
      net674, net673, net672, net671, net670, net669, net668, net667, net666, 
      net665, net664, net663, net662, net661, net660, net659, net658, net657, 
      net656, net655, net654, net653, net652, net651, net650, net649, net648, 
      net647, net646, net645, net644, net643, net642, net641, net640, net639, 
      net638, net637, net636, net635, net634, net633, net632, net631, net630, 
      net629, net628, net627, net626, net625, net624, net623, net622, net621, 
      net620, net619, net618, net617, net616, net615, net614, net613, net612, 
      net611, net610, net609, net608, net607, net606, net605, net604, net603, 
      net602, net601, net600, net599, net598, net597, net596, net595, net594, 
      net593, net592, net591, net590, net589, net588, net587, net586, n168, 
      n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, 
      n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, 
      n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, 
      n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, 
      n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, 
      n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, 
      n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, 
      n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, 
      n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, 
      n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288, 
      n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, net43112, 
      net43113, net43114 : std_logic;

begin
   
   X_Logic1_port <= '1';
   X_Logic0_port <= '0';
   n1 <= '0';
   n2 <= '0';
   npc2_reg_0_inst : DFFR_X1 port map( D => n296, CK => Clk, RN => Rst, Q => 
                           npc2_0_port, QN => net586);
   PC_reg_31_inst : DFFR_X1 port map( D => n295, CK => Clk, RN => Rst, Q => 
                           PC_31_port, QN => net681);
   out_NPC_reg_31_inst : DFFR_X1 port map( D => n294, CK => Clk, RN => Rst, Q 
                           => out_NPC_31_port, QN => net649);
   npc2_reg_31_inst : DFFR_X1 port map( D => n293, CK => Clk, RN => Rst, Q => 
                           npc2_31_port, QN => net617);
   out_NPC_reg_0_inst : DFFR_X1 port map( D => n292, CK => Clk, RN => Rst, Q =>
                           out_NPC_0_port, QN => net618);
   out_NPC_reg_1_inst : DFFR_X1 port map( D => n291, CK => Clk, RN => Rst, Q =>
                           out_NPC_1_port, QN => net619);
   npc2_reg_1_inst : DFFR_X1 port map( D => n290, CK => Clk, RN => Rst, Q => 
                           npc2_1_port, QN => net587);
   out_NPC_reg_2_inst : DFFR_X1 port map( D => n289, CK => Clk, RN => Rst, Q =>
                           out_NPC_2_port, QN => net620);
   npc2_reg_2_inst : DFFR_X1 port map( D => n288, CK => Clk, RN => Rst, Q => 
                           npc2_2_port, QN => net588);
   out_NPC_reg_3_inst : DFFR_X1 port map( D => n287, CK => Clk, RN => Rst, Q =>
                           out_NPC_3_port, QN => net621);
   npc2_reg_3_inst : DFFR_X1 port map( D => n286, CK => Clk, RN => Rst, Q => 
                           npc2_3_port, QN => net589);
   out_NPC_reg_4_inst : DFFR_X1 port map( D => n285, CK => Clk, RN => Rst, Q =>
                           out_NPC_4_port, QN => net622);
   npc2_reg_4_inst : DFFR_X1 port map( D => n284, CK => Clk, RN => Rst, Q => 
                           npc2_4_port, QN => net590);
   out_NPC_reg_5_inst : DFFR_X1 port map( D => n283, CK => Clk, RN => Rst, Q =>
                           out_NPC_5_port, QN => net623);
   npc2_reg_5_inst : DFFR_X1 port map( D => n282, CK => Clk, RN => Rst, Q => 
                           npc2_5_port, QN => net591);
   out_NPC_reg_6_inst : DFFR_X1 port map( D => n281, CK => Clk, RN => Rst, Q =>
                           out_NPC_6_port, QN => net624);
   npc2_reg_6_inst : DFFR_X1 port map( D => n280, CK => Clk, RN => Rst, Q => 
                           npc2_6_port, QN => net592);
   out_NPC_reg_7_inst : DFFR_X1 port map( D => n279, CK => Clk, RN => Rst, Q =>
                           out_NPC_7_port, QN => net625);
   npc2_reg_7_inst : DFFR_X1 port map( D => n278, CK => Clk, RN => Rst, Q => 
                           npc2_7_port, QN => net593);
   out_NPC_reg_8_inst : DFFR_X1 port map( D => n277, CK => Clk, RN => Rst, Q =>
                           out_NPC_8_port, QN => net626);
   npc2_reg_8_inst : DFFR_X1 port map( D => n276, CK => Clk, RN => Rst, Q => 
                           npc2_8_port, QN => net594);
   out_NPC_reg_9_inst : DFFR_X1 port map( D => n275, CK => Clk, RN => Rst, Q =>
                           out_NPC_9_port, QN => net627);
   npc2_reg_9_inst : DFFR_X1 port map( D => n274, CK => Clk, RN => Rst, Q => 
                           npc2_9_port, QN => net595);
   out_NPC_reg_10_inst : DFFR_X1 port map( D => n273, CK => Clk, RN => Rst, Q 
                           => out_NPC_10_port, QN => net628);
   npc2_reg_10_inst : DFFR_X1 port map( D => n272, CK => Clk, RN => Rst, Q => 
                           npc2_10_port, QN => net596);
   out_NPC_reg_11_inst : DFFR_X1 port map( D => n271, CK => Clk, RN => Rst, Q 
                           => out_NPC_11_port, QN => net629);
   npc2_reg_11_inst : DFFR_X1 port map( D => n270, CK => Clk, RN => Rst, Q => 
                           npc2_11_port, QN => net597);
   out_NPC_reg_12_inst : DFFR_X1 port map( D => n269, CK => Clk, RN => Rst, Q 
                           => out_NPC_12_port, QN => net630);
   npc2_reg_12_inst : DFFR_X1 port map( D => n268, CK => Clk, RN => Rst, Q => 
                           npc2_12_port, QN => net598);
   out_NPC_reg_13_inst : DFFR_X1 port map( D => n267, CK => Clk, RN => Rst, Q 
                           => out_NPC_13_port, QN => net631);
   npc2_reg_13_inst : DFFR_X1 port map( D => n266, CK => Clk, RN => Rst, Q => 
                           npc2_13_port, QN => net599);
   out_NPC_reg_14_inst : DFFR_X1 port map( D => n265, CK => Clk, RN => Rst, Q 
                           => out_NPC_14_port, QN => net632);
   npc2_reg_14_inst : DFFR_X1 port map( D => n264, CK => Clk, RN => Rst, Q => 
                           npc2_14_port, QN => net600);
   out_NPC_reg_15_inst : DFFR_X1 port map( D => n263, CK => Clk, RN => Rst, Q 
                           => out_NPC_15_port, QN => net633);
   npc2_reg_15_inst : DFFR_X1 port map( D => n262, CK => Clk, RN => Rst, Q => 
                           npc2_15_port, QN => net601);
   out_NPC_reg_16_inst : DFFR_X1 port map( D => n261, CK => Clk, RN => Rst, Q 
                           => out_NPC_16_port, QN => net634);
   npc2_reg_16_inst : DFFR_X1 port map( D => n260, CK => Clk, RN => Rst, Q => 
                           npc2_16_port, QN => net602);
   out_NPC_reg_17_inst : DFFR_X1 port map( D => n259, CK => Clk, RN => Rst, Q 
                           => out_NPC_17_port, QN => net635);
   npc2_reg_17_inst : DFFR_X1 port map( D => n258, CK => Clk, RN => Rst, Q => 
                           npc2_17_port, QN => net603);
   out_NPC_reg_18_inst : DFFR_X1 port map( D => n257, CK => Clk, RN => Rst, Q 
                           => out_NPC_18_port, QN => net636);
   npc2_reg_18_inst : DFFR_X1 port map( D => n256, CK => Clk, RN => Rst, Q => 
                           npc2_18_port, QN => net604);
   out_NPC_reg_19_inst : DFFR_X1 port map( D => n255, CK => Clk, RN => Rst, Q 
                           => out_NPC_19_port, QN => net637);
   npc2_reg_19_inst : DFFR_X1 port map( D => n254, CK => Clk, RN => Rst, Q => 
                           npc2_19_port, QN => net605);
   out_NPC_reg_20_inst : DFFR_X1 port map( D => n253, CK => Clk, RN => Rst, Q 
                           => out_NPC_20_port, QN => net638);
   npc2_reg_20_inst : DFFR_X1 port map( D => n252, CK => Clk, RN => Rst, Q => 
                           npc2_20_port, QN => net606);
   out_NPC_reg_21_inst : DFFR_X1 port map( D => n251, CK => Clk, RN => Rst, Q 
                           => out_NPC_21_port, QN => net639);
   npc2_reg_21_inst : DFFR_X1 port map( D => n250, CK => Clk, RN => Rst, Q => 
                           npc2_21_port, QN => net607);
   out_NPC_reg_22_inst : DFFR_X1 port map( D => n249, CK => Clk, RN => Rst, Q 
                           => out_NPC_22_port, QN => net640);
   npc2_reg_22_inst : DFFR_X1 port map( D => n248, CK => Clk, RN => Rst, Q => 
                           npc2_22_port, QN => net608);
   out_NPC_reg_23_inst : DFFR_X1 port map( D => n247, CK => Clk, RN => Rst, Q 
                           => out_NPC_23_port, QN => net641);
   npc2_reg_23_inst : DFFR_X1 port map( D => n246, CK => Clk, RN => Rst, Q => 
                           npc2_23_port, QN => net609);
   out_NPC_reg_24_inst : DFFR_X1 port map( D => n245, CK => Clk, RN => Rst, Q 
                           => out_NPC_24_port, QN => net642);
   npc2_reg_24_inst : DFFR_X1 port map( D => n244, CK => Clk, RN => Rst, Q => 
                           npc2_24_port, QN => net610);
   out_NPC_reg_25_inst : DFFR_X1 port map( D => n243, CK => Clk, RN => Rst, Q 
                           => out_NPC_25_port, QN => net643);
   npc2_reg_25_inst : DFFR_X1 port map( D => n242, CK => Clk, RN => Rst, Q => 
                           npc2_25_port, QN => net611);
   out_NPC_reg_26_inst : DFFR_X1 port map( D => n241, CK => Clk, RN => Rst, Q 
                           => out_NPC_26_port, QN => net644);
   npc2_reg_26_inst : DFFR_X1 port map( D => n240, CK => Clk, RN => Rst, Q => 
                           npc2_26_port, QN => net612);
   out_NPC_reg_27_inst : DFFR_X1 port map( D => n239, CK => Clk, RN => Rst, Q 
                           => out_NPC_27_port, QN => net645);
   npc2_reg_27_inst : DFFR_X1 port map( D => n238, CK => Clk, RN => Rst, Q => 
                           npc2_27_port, QN => net613);
   out_NPC_reg_28_inst : DFFR_X1 port map( D => n237, CK => Clk, RN => Rst, Q 
                           => out_NPC_28_port, QN => net646);
   npc2_reg_28_inst : DFFR_X1 port map( D => n236, CK => Clk, RN => Rst, Q => 
                           npc2_28_port, QN => net614);
   out_NPC_reg_29_inst : DFFR_X1 port map( D => n235, CK => Clk, RN => Rst, Q 
                           => out_NPC_29_port, QN => net647);
   npc2_reg_29_inst : DFFR_X1 port map( D => n234, CK => Clk, RN => Rst, Q => 
                           npc2_29_port, QN => net615);
   out_NPC_reg_30_inst : DFFR_X1 port map( D => n233, CK => Clk, RN => Rst, Q 
                           => out_NPC_30_port, QN => net648);
   npc2_reg_30_inst : DFFR_X1 port map( D => n232, CK => Clk, RN => Rst, Q => 
                           npc2_30_port, QN => net616);
   PC_reg_0_inst : DFFR_X1 port map( D => n231, CK => Clk, RN => Rst, Q => 
                           PC_0_port, QN => net650);
   PC_reg_1_inst : DFFR_X1 port map( D => n230, CK => Clk, RN => Rst, Q => 
                           PC_1_port, QN => net651);
   PC_reg_2_inst : DFFR_X1 port map( D => n229, CK => Clk, RN => Rst, Q => 
                           PC_2_port, QN => net652);
   PC_reg_3_inst : DFFR_X1 port map( D => n228, CK => Clk, RN => Rst, Q => 
                           PC_3_port, QN => net653);
   PC_reg_4_inst : DFFR_X1 port map( D => n227, CK => Clk, RN => Rst, Q => 
                           PC_4_port, QN => net654);
   PC_reg_5_inst : DFFR_X1 port map( D => n226, CK => Clk, RN => Rst, Q => 
                           PC_5_port, QN => net655);
   PC_reg_6_inst : DFFR_X1 port map( D => n225, CK => Clk, RN => Rst, Q => 
                           PC_6_port, QN => net656);
   PC_reg_7_inst : DFFR_X1 port map( D => n224, CK => Clk, RN => Rst, Q => 
                           PC_7_port, QN => net657);
   PC_reg_8_inst : DFFR_X1 port map( D => n223, CK => Clk, RN => Rst, Q => 
                           PC_8_port, QN => net658);
   PC_reg_9_inst : DFFR_X1 port map( D => n222, CK => Clk, RN => Rst, Q => 
                           PC_9_port, QN => net659);
   PC_reg_10_inst : DFFR_X1 port map( D => n221, CK => Clk, RN => Rst, Q => 
                           PC_10_port, QN => net660);
   PC_reg_11_inst : DFFR_X1 port map( D => n220, CK => Clk, RN => Rst, Q => 
                           PC_11_port, QN => net661);
   PC_reg_12_inst : DFFR_X1 port map( D => n219, CK => Clk, RN => Rst, Q => 
                           PC_12_port, QN => net662);
   PC_reg_13_inst : DFFR_X1 port map( D => n218, CK => Clk, RN => Rst, Q => 
                           PC_13_port, QN => net663);
   PC_reg_14_inst : DFFR_X1 port map( D => n217, CK => Clk, RN => Rst, Q => 
                           PC_14_port, QN => net664);
   PC_reg_15_inst : DFFR_X1 port map( D => n216, CK => Clk, RN => Rst, Q => 
                           PC_15_port, QN => net665);
   PC_reg_16_inst : DFFR_X1 port map( D => n215, CK => Clk, RN => Rst, Q => 
                           PC_16_port, QN => net666);
   PC_reg_17_inst : DFFR_X1 port map( D => n214, CK => Clk, RN => Rst, Q => 
                           PC_17_port, QN => net667);
   PC_reg_18_inst : DFFR_X1 port map( D => n213, CK => Clk, RN => Rst, Q => 
                           PC_18_port, QN => net668);
   PC_reg_19_inst : DFFR_X1 port map( D => n212, CK => Clk, RN => Rst, Q => 
                           PC_19_port, QN => net669);
   PC_reg_20_inst : DFFR_X1 port map( D => n211, CK => Clk, RN => Rst, Q => 
                           PC_20_port, QN => net670);
   PC_reg_21_inst : DFFR_X1 port map( D => n210, CK => Clk, RN => Rst, Q => 
                           PC_21_port, QN => net671);
   PC_reg_22_inst : DFFR_X1 port map( D => n209, CK => Clk, RN => Rst, Q => 
                           PC_22_port, QN => net672);
   PC_reg_23_inst : DFFR_X1 port map( D => n208, CK => Clk, RN => Rst, Q => 
                           PC_23_port, QN => net673);
   PC_reg_24_inst : DFFR_X1 port map( D => n207, CK => Clk, RN => Rst, Q => 
                           PC_24_port, QN => net674);
   PC_reg_25_inst : DFFR_X1 port map( D => n206, CK => Clk, RN => Rst, Q => 
                           PC_25_port, QN => net675);
   PC_reg_26_inst : DFFR_X1 port map( D => n205, CK => Clk, RN => Rst, Q => 
                           PC_26_port, QN => net676);
   PC_reg_27_inst : DFFR_X1 port map( D => n204, CK => Clk, RN => Rst, Q => 
                           PC_27_port, QN => net677);
   PC_reg_28_inst : DFFR_X1 port map( D => n203, CK => Clk, RN => Rst, Q => 
                           PC_28_port, QN => net678);
   PC_reg_29_inst : DFFR_X1 port map( D => n202, CK => Clk, RN => Rst, Q => 
                           PC_29_port, QN => net679);
   PC_reg_30_inst : DFFR_X1 port map( D => n201, CK => Clk, RN => Rst, Q => 
                           PC_30_port, QN => net680);
   IR_reg_7_inst : DFFR_X1 port map( D => n200, CK => Clk, RN => n168, Q => 
                           IR_7_port, QN => net689);
   IR_reg_5_inst : DFFR_X1 port map( D => n199, CK => Clk, RN => n168, Q => 
                           IR_5_port, QN => net687);
   IR_reg_3_inst : DFFR_X1 port map( D => n198, CK => Clk, RN => n168, Q => 
                           IR_3_port, QN => net685);
   IR_reg_31_inst : DFFR_X1 port map( D => n197, CK => Clk, RN => n168, Q => 
                           IR_31_port, QN => net713);
   IR_reg_29_inst : DFFR_X1 port map( D => n196, CK => Clk, RN => n168, Q => 
                           IR_29_port, QN => net711);
   IR_reg_1_inst : DFFR_X1 port map( D => n195, CK => Clk, RN => n168, Q => 
                           IR_1_port, QN => net683);
   IR_reg_26_inst : DFFR_X1 port map( D => n194, CK => Clk, RN => n168, Q => 
                           IR_26_port, QN => net708);
   IR_reg_24_inst : DFFR_X1 port map( D => n193, CK => Clk, RN => n168, Q => 
                           IR_24_port, QN => net706);
   IR_reg_22_inst : DFFR_X1 port map( D => n192, CK => Clk, RN => n168, Q => 
                           IR_22_port, QN => net704);
   IR_reg_20_inst : DFFR_X1 port map( D => n191, CK => Clk, RN => n168, Q => 
                           IR_20_port, QN => net702);
   IR_reg_18_inst : DFFR_X1 port map( D => n190, CK => Clk, RN => n168, Q => 
                           IR_18_port, QN => net700);
   IR_reg_17_inst : DFFR_X1 port map( D => n189, CK => Clk, RN => n168, Q => 
                           IR_17_port, QN => net699);
   IR_reg_15_inst : DFFR_X1 port map( D => n188, CK => Clk, RN => n168, Q => 
                           IR_15_port, QN => net697);
   IR_reg_13_inst : DFFR_X1 port map( D => n187, CK => Clk, RN => n168, Q => 
                           IR_13_port, QN => net695);
   IR_reg_11_inst : DFFR_X1 port map( D => n186, CK => Clk, RN => n168, Q => 
                           IR_11_port, QN => net693);
   IR_reg_9_inst : DFFR_X1 port map( D => n185, CK => Clk, RN => n168, Q => 
                           IR_9_port, QN => net691);
   IR_reg_8_inst : DFFR_X1 port map( D => n184, CK => Clk, RN => n168, Q => 
                           IR_8_port, QN => net690);
   IR_reg_10_inst : DFFR_X1 port map( D => n183, CK => Clk, RN => n168, Q => 
                           IR_10_port, QN => net692);
   IR_reg_12_inst : DFFR_X1 port map( D => n182, CK => Clk, RN => n168, Q => 
                           IR_12_port, QN => net694);
   IR_reg_14_inst : DFFR_X1 port map( D => n181, CK => Clk, RN => n168, Q => 
                           IR_14_port, QN => net696);
   IR_reg_16_inst : DFFR_X1 port map( D => n180, CK => Clk, RN => n168, Q => 
                           IR_16_port, QN => net698);
   IR_reg_0_inst : DFFR_X1 port map( D => n179, CK => Clk, RN => n168, Q => 
                           IR_0_port, QN => net682);
   IR_reg_19_inst : DFFR_X1 port map( D => n178, CK => Clk, RN => n168, Q => 
                           IR_19_port, QN => net701);
   IR_reg_21_inst : DFFR_X1 port map( D => n177, CK => Clk, RN => n168, Q => 
                           IR_21_port, QN => net703);
   IR_reg_23_inst : DFFR_X1 port map( D => n176, CK => Clk, RN => n168, Q => 
                           IR_23_port, QN => net705);
   IR_reg_25_inst : DFFR_X1 port map( D => n175, CK => Clk, RN => n168, Q => 
                           IR_25_port, QN => net707);
   IR_reg_27_inst : DFFR_X1 port map( D => n174, CK => Clk, RN => n168, Q => 
                           IR_27_port, QN => net709);
   IR_reg_28_inst : DFFR_X1 port map( D => n173, CK => Clk, RN => n168, Q => 
                           IR_28_port, QN => net710);
   IR_reg_30_inst : DFFR_X1 port map( D => n172, CK => Clk, RN => n168, Q => 
                           IR_30_port, QN => net712);
   IR_reg_2_inst : DFFR_X1 port map( D => n171, CK => Clk, RN => n168, Q => 
                           IR_2_port, QN => net684);
   IR_reg_4_inst : DFFR_X1 port map( D => n170, CK => Clk, RN => n168, Q => 
                           IR_4_port, QN => net686);
   IR_reg_6_inst : DFFR_X1 port map( D => n169, CK => Clk, RN => n168, Q => 
                           IR_6_port, QN => net688);
   DP_I : datapath_reg_size32 port map( clk => Clk, rst => Rst, flush => 
                           jump_verified, RF1 => rd1_i, RF2 => rd2_i, WF1 => 
                           wr_i, EN_regA => RegA_LATCH_EN_i, EN_regB => 
                           RegB_LATCH_EN_i, EN_regIMM => RegIMM_LATCH_EN_i, 
                           EN_regALUOP => RegAluOpCodeGen_EN_i, EN_regRD1 => 
                           en_RD1_i, EN_regNPC2 => NPC2_LATCH_EN_i, S1 => 
                           MUXA_SEL_i, S2 => MUXB_SEL_i, EN_regRET => 
                           RETURN_REG_EN_i, EN_regOUTALU => ALU_OUTREG_EN_i, 
                           EN_regB2 => B2_EN_i, EN_regRD2 => en_RD2_i, 
                           EN_regALU2 => Alu_outreg2_en_i, EN_regLMD => 
                           LMD_LATCH_EN_i, EN_regRD3 => en_RD3_i, Sel_ret_alu 
                           => sel_alu_ret_i, Sel_alu_lmd => WB_MUX_SEL_i, 
                           sel_31_rd => wb_mux_add_sel_i, NPC(31) => 
                           out_NPC_31_port, NPC(30) => out_NPC_30_port, NPC(29)
                           => out_NPC_29_port, NPC(28) => out_NPC_28_port, 
                           NPC(27) => out_NPC_27_port, NPC(26) => 
                           out_NPC_26_port, NPC(25) => out_NPC_25_port, NPC(24)
                           => out_NPC_24_port, NPC(23) => out_NPC_23_port, 
                           NPC(22) => out_NPC_22_port, NPC(21) => 
                           out_NPC_21_port, NPC(20) => out_NPC_20_port, NPC(19)
                           => out_NPC_19_port, NPC(18) => out_NPC_18_port, 
                           NPC(17) => out_NPC_17_port, NPC(16) => 
                           out_NPC_16_port, NPC(15) => out_NPC_15_port, NPC(14)
                           => out_NPC_14_port, NPC(13) => out_NPC_13_port, 
                           NPC(12) => out_NPC_12_port, NPC(11) => 
                           out_NPC_11_port, NPC(10) => out_NPC_10_port, NPC(9) 
                           => out_NPC_9_port, NPC(8) => out_NPC_8_port, NPC(7) 
                           => out_NPC_7_port, NPC(6) => out_NPC_6_port, NPC(5) 
                           => out_NPC_5_port, NPC(4) => out_NPC_4_port, NPC(3) 
                           => out_NPC_3_port, NPC(2) => out_NPC_2_port, NPC(1) 
                           => out_NPC_1_port, NPC(0) => out_NPC_0_port, 
                           IR_dp(31) => IR_31_port, IR_dp(30) => IR_30_port, 
                           IR_dp(29) => IR_29_port, IR_dp(28) => IR_28_port, 
                           IR_dp(27) => IR_27_port, IR_dp(26) => IR_26_port, 
                           IR_dp(25) => IR_25_port, IR_dp(24) => IR_24_port, 
                           IR_dp(23) => IR_23_port, IR_dp(22) => IR_22_port, 
                           IR_dp(21) => IR_21_port, IR_dp(20) => IR_20_port, 
                           IR_dp(19) => IR_19_port, IR_dp(18) => IR_18_port, 
                           IR_dp(17) => IR_17_port, IR_dp(16) => IR_16_port, 
                           IR_dp(15) => IR_15_port, IR_dp(14) => IR_14_port, 
                           IR_dp(13) => IR_13_port, IR_dp(12) => IR_12_port, 
                           IR_dp(11) => IR_11_port, IR_dp(10) => IR_10_port, 
                           IR_dp(9) => IR_9_port, IR_dp(8) => IR_8_port, 
                           IR_dp(7) => IR_7_port, IR_dp(6) => IR_6_port, 
                           IR_dp(5) => IR_5_port, IR_dp(4) => IR_4_port, 
                           IR_dp(3) => IR_3_port, IR_dp(2) => IR_2_port, 
                           IR_dp(1) => IR_1_port, IR_dp(0) => IR_0_port, 
                           OUT_DP(31) => net714, OUT_DP(30) => net715, 
                           OUT_DP(29) => net716, OUT_DP(28) => net717, 
                           OUT_DP(27) => net718, OUT_DP(26) => net719, 
                           OUT_DP(25) => net720, OUT_DP(24) => net721, 
                           OUT_DP(23) => net722, OUT_DP(22) => net723, 
                           OUT_DP(21) => net724, OUT_DP(20) => net725, 
                           OUT_DP(19) => net726, OUT_DP(18) => net727, 
                           OUT_DP(17) => net728, OUT_DP(16) => net729, 
                           OUT_DP(15) => net730, OUT_DP(14) => net731, 
                           OUT_DP(13) => net732, OUT_DP(12) => net733, 
                           OUT_DP(11) => net734, OUT_DP(10) => net735, 
                           OUT_DP(9) => net736, OUT_DP(8) => net737, OUT_DP(7) 
                           => net738, OUT_DP(6) => net739, OUT_DP(5) => net740,
                           OUT_DP(4) => net741, OUT_DP(3) => net742, OUT_DP(2) 
                           => net743, OUT_DP(1) => net744, OUT_DP(0) => net745,
                           comp_branch_i => comp_branch_dp, 
                           immediate_branch(31) => immediate_31_port, 
                           immediate_branch(30) => immediate_30_port, 
                           immediate_branch(29) => immediate_29_port, 
                           immediate_branch(28) => immediate_28_port, 
                           immediate_branch(27) => immediate_27_port, 
                           immediate_branch(26) => immediate_26_port, 
                           immediate_branch(25) => immediate_25_port, 
                           immediate_branch(24) => immediate_24_port, 
                           immediate_branch(23) => immediate_23_port, 
                           immediate_branch(22) => immediate_22_port, 
                           immediate_branch(21) => immediate_21_port, 
                           immediate_branch(20) => immediate_20_port, 
                           immediate_branch(19) => immediate_19_port, 
                           immediate_branch(18) => immediate_18_port, 
                           immediate_branch(17) => immediate_17_port, 
                           immediate_branch(16) => immediate_16_port, 
                           immediate_branch(15) => immediate_15_port, 
                           immediate_branch(14) => immediate_14_port, 
                           immediate_branch(13) => immediate_13_port, 
                           immediate_branch(12) => immediate_12_port, 
                           immediate_branch(11) => immediate_11_port, 
                           immediate_branch(10) => immediate_10_port, 
                           immediate_branch(9) => immediate_9_port, 
                           immediate_branch(8) => immediate_8_port, 
                           immediate_branch(7) => immediate_7_port, 
                           immediate_branch(6) => immediate_6_port, 
                           immediate_branch(5) => immediate_5_port, 
                           immediate_branch(4) => immediate_4_port, 
                           immediate_branch(3) => immediate_3_port, 
                           immediate_branch(2) => immediate_2_port, 
                           immediate_branch(1) => immediate_1_port, 
                           immediate_branch(0) => immediate_0_port, ADD_mem(31)
                           => dram_ADD(31), ADD_mem(30) => dram_ADD(30), 
                           ADD_mem(29) => dram_ADD(29), ADD_mem(28) => 
                           dram_ADD(28), ADD_mem(27) => dram_ADD(27), 
                           ADD_mem(26) => dram_ADD(26), ADD_mem(25) => 
                           dram_ADD(25), ADD_mem(24) => dram_ADD(24), 
                           ADD_mem(23) => dram_ADD(23), ADD_mem(22) => 
                           dram_ADD(22), ADD_mem(21) => dram_ADD(21), 
                           ADD_mem(20) => dram_ADD(20), ADD_mem(19) => 
                           dram_ADD(19), ADD_mem(18) => dram_ADD(18), 
                           ADD_mem(17) => dram_ADD(17), ADD_mem(16) => 
                           dram_ADD(16), ADD_mem(15) => dram_ADD(15), 
                           ADD_mem(14) => dram_ADD(14), ADD_mem(13) => 
                           dram_ADD(13), ADD_mem(12) => dram_ADD(12), 
                           ADD_mem(11) => dram_ADD(11), ADD_mem(10) => 
                           dram_ADD(10), ADD_mem(9) => dram_ADD(9), ADD_mem(8) 
                           => dram_ADD(8), ADD_mem(7) => dram_ADD(7), 
                           ADD_mem(6) => dram_ADD(6), ADD_mem(5) => dram_ADD(5)
                           , ADD_mem(4) => dram_ADD(4), ADD_mem(3) => 
                           dram_ADD(3), ADD_mem(2) => dram_ADD(2), ADD_mem(1) 
                           => dram_ADD(1), ADD_mem(0) => dram_ADD(0), 
                           DIN_mem(31) => dram_DIN(31), DIN_mem(30) => 
                           dram_DIN(30), DIN_mem(29) => dram_DIN(29), 
                           DIN_mem(28) => dram_DIN(28), DIN_mem(27) => 
                           dram_DIN(27), DIN_mem(26) => dram_DIN(26), 
                           DIN_mem(25) => dram_DIN(25), DIN_mem(24) => 
                           dram_DIN(24), DIN_mem(23) => dram_DIN(23), 
                           DIN_mem(22) => dram_DIN(22), DIN_mem(21) => 
                           dram_DIN(21), DIN_mem(20) => dram_DIN(20), 
                           DIN_mem(19) => dram_DIN(19), DIN_mem(18) => 
                           dram_DIN(18), DIN_mem(17) => dram_DIN(17), 
                           DIN_mem(16) => dram_DIN(16), DIN_mem(15) => 
                           dram_DIN(15), DIN_mem(14) => dram_DIN(14), 
                           DIN_mem(13) => dram_DIN(13), DIN_mem(12) => 
                           dram_DIN(12), DIN_mem(11) => dram_DIN(11), 
                           DIN_mem(10) => dram_DIN(10), DIN_mem(9) => 
                           dram_DIN(9), DIN_mem(8) => dram_DIN(8), DIN_mem(7) 
                           => dram_DIN(7), DIN_mem(6) => dram_DIN(6), 
                           DIN_mem(5) => dram_DIN(5), DIN_mem(4) => dram_DIN(4)
                           , DIN_mem(3) => dram_DIN(3), DIN_mem(2) => 
                           dram_DIN(2), DIN_mem(1) => dram_DIN(1), DIN_mem(0) 
                           => dram_DIN(0), DOUT_mem(31) => dram_DOUT(31), 
                           DOUT_mem(30) => dram_DOUT(30), DOUT_mem(29) => 
                           dram_DOUT(29), DOUT_mem(28) => dram_DOUT(28), 
                           DOUT_mem(27) => dram_DOUT(27), DOUT_mem(26) => 
                           dram_DOUT(26), DOUT_mem(25) => dram_DOUT(25), 
                           DOUT_mem(24) => dram_DOUT(24), DOUT_mem(23) => 
                           dram_DOUT(23), DOUT_mem(22) => dram_DOUT(22), 
                           DOUT_mem(21) => dram_DOUT(21), DOUT_mem(20) => 
                           dram_DOUT(20), DOUT_mem(19) => dram_DOUT(19), 
                           DOUT_mem(18) => dram_DOUT(18), DOUT_mem(17) => 
                           dram_DOUT(17), DOUT_mem(16) => dram_DOUT(16), 
                           DOUT_mem(15) => dram_DOUT(15), DOUT_mem(14) => 
                           dram_DOUT(14), DOUT_mem(13) => dram_DOUT(13), 
                           DOUT_mem(12) => dram_DOUT(12), DOUT_mem(11) => 
                           dram_DOUT(11), DOUT_mem(10) => dram_DOUT(10), 
                           DOUT_mem(9) => dram_DOUT(9), DOUT_mem(8) => 
                           dram_DOUT(8), DOUT_mem(7) => dram_DOUT(7), 
                           DOUT_mem(6) => dram_DOUT(6), DOUT_mem(5) => 
                           dram_DOUT(5), DOUT_mem(4) => dram_DOUT(4), 
                           DOUT_mem(3) => dram_DOUT(3), DOUT_mem(2) => 
                           dram_DOUT(2), DOUT_mem(1) => dram_DOUT(1), 
                           DOUT_mem(0) => dram_DOUT(0));
   mux_pc : mux21_N32_0 port map( A(31) => in_NPC_31_port, A(30) => 
                           in_NPC_30_port, A(29) => in_NPC_29_port, A(28) => 
                           in_NPC_28_port, A(27) => in_NPC_27_port, A(26) => 
                           in_NPC_26_port, A(25) => in_NPC_25_port, A(24) => 
                           in_NPC_24_port, A(23) => in_NPC_23_port, A(22) => 
                           in_NPC_22_port, A(21) => in_NPC_21_port, A(20) => 
                           in_NPC_20_port, A(19) => in_NPC_19_port, A(18) => 
                           in_NPC_18_port, A(17) => in_NPC_17_port, A(16) => 
                           in_NPC_16_port, A(15) => in_NPC_15_port, A(14) => 
                           in_NPC_14_port, A(13) => in_NPC_13_port, A(12) => 
                           in_NPC_12_port, A(11) => in_NPC_11_port, A(10) => 
                           in_NPC_10_port, A(9) => in_NPC_9_port, A(8) => 
                           in_NPC_8_port, A(7) => in_NPC_7_port, A(6) => 
                           in_NPC_6_port, A(5) => in_NPC_5_port, A(4) => 
                           in_NPC_4_port, A(3) => in_NPC_3_port, A(2) => 
                           in_NPC_2_port, A(1) => in_NPC_1_port, A(0) => 
                           in_NPC_0_port, B(31) => pc_jump_31_port, B(30) => 
                           pc_jump_30_port, B(29) => pc_jump_29_port, B(28) => 
                           pc_jump_28_port, B(27) => pc_jump_27_port, B(26) => 
                           pc_jump_26_port, B(25) => pc_jump_25_port, B(24) => 
                           pc_jump_24_port, B(23) => pc_jump_23_port, B(22) => 
                           pc_jump_22_port, B(21) => pc_jump_21_port, B(20) => 
                           pc_jump_20_port, B(19) => pc_jump_19_port, B(18) => 
                           pc_jump_18_port, B(17) => pc_jump_17_port, B(16) => 
                           pc_jump_16_port, B(15) => pc_jump_15_port, B(14) => 
                           pc_jump_14_port, B(13) => pc_jump_13_port, B(12) => 
                           pc_jump_12_port, B(11) => pc_jump_11_port, B(10) => 
                           pc_jump_10_port, B(9) => pc_jump_9_port, B(8) => 
                           pc_jump_8_port, B(7) => pc_jump_7_port, B(6) => 
                           pc_jump_6_port, B(5) => pc_jump_5_port, B(4) => 
                           pc_jump_4_port, B(3) => pc_jump_3_port, B(2) => 
                           pc_jump_2_port, B(1) => pc_jump_1_port, B(0) => 
                           pc_jump_0_port, SEL => jump_verified, Y(31) => 
                           PC_BUS_31_port, Y(30) => PC_BUS_30_port, Y(29) => 
                           PC_BUS_29_port, Y(28) => PC_BUS_28_port, Y(27) => 
                           PC_BUS_27_port, Y(26) => PC_BUS_26_port, Y(25) => 
                           PC_BUS_25_port, Y(24) => PC_BUS_24_port, Y(23) => 
                           PC_BUS_23_port, Y(22) => PC_BUS_22_port, Y(21) => 
                           PC_BUS_21_port, Y(20) => PC_BUS_20_port, Y(19) => 
                           PC_BUS_19_port, Y(18) => PC_BUS_18_port, Y(17) => 
                           PC_BUS_17_port, Y(16) => PC_BUS_16_port, Y(15) => 
                           PC_BUS_15_port, Y(14) => PC_BUS_14_port, Y(13) => 
                           PC_BUS_13_port, Y(12) => PC_BUS_12_port, Y(11) => 
                           PC_BUS_11_port, Y(10) => PC_BUS_10_port, Y(9) => 
                           PC_BUS_9_port, Y(8) => PC_BUS_8_port, Y(7) => 
                           PC_BUS_7_port, Y(6) => PC_BUS_6_port, Y(5) => 
                           PC_BUS_5_port, Y(4) => PC_BUS_4_port, Y(3) => 
                           PC_BUS_3_port, Y(2) => PC_BUS_2_port, Y(1) => 
                           PC_BUS_1_port, Y(0) => PC_BUS_0_port);
   CU_I : 
                           CU_HDW_MICROCODE_MEM_SIZE10_FUNC_SIZE11_OP_CODE_SIZE6_IR_SIZE32_CW_SIZE21 
                           port map( Clk => Clk, Rst => Rst, IR_IN(31) => 
                           iram_Dout(31), IR_IN(30) => iram_Dout(30), IR_IN(29)
                           => iram_Dout(29), IR_IN(28) => iram_Dout(28), 
                           IR_IN(27) => iram_Dout(27), IR_IN(26) => 
                           iram_Dout(26), IR_IN(25) => iram_Dout(25), IR_IN(24)
                           => iram_Dout(24), IR_IN(23) => iram_Dout(23), 
                           IR_IN(22) => iram_Dout(22), IR_IN(21) => 
                           iram_Dout(21), IR_IN(20) => iram_Dout(20), IR_IN(19)
                           => iram_Dout(19), IR_IN(18) => iram_Dout(18), 
                           IR_IN(17) => iram_Dout(17), IR_IN(16) => 
                           iram_Dout(16), IR_IN(15) => iram_Dout(15), IR_IN(14)
                           => iram_Dout(14), IR_IN(13) => iram_Dout(13), 
                           IR_IN(12) => iram_Dout(12), IR_IN(11) => 
                           iram_Dout(11), IR_IN(10) => iram_Dout(10), IR_IN(9) 
                           => iram_Dout(9), IR_IN(8) => iram_Dout(8), IR_IN(7) 
                           => iram_Dout(7), IR_IN(6) => iram_Dout(6), IR_IN(5) 
                           => iram_Dout(5), IR_IN(4) => iram_Dout(4), IR_IN(3) 
                           => iram_Dout(3), IR_IN(2) => iram_Dout(2), IR_IN(1) 
                           => iram_Dout(1), IR_IN(0) => iram_Dout(0), flush => 
                           jump_verified, IR_LATCH_EN => net43114, 
                           NPC1_LATCH_EN => NPC1_LATCH_EN_i, NPC2_LATCH_EN => 
                           NPC2_LATCH_EN_i, RegA_LATCH_EN => RegA_LATCH_EN_i, 
                           RegB_LATCH_EN => RegB_LATCH_EN_i, RegAluOpCodeGen_EN
                           => RegAluOpCodeGen_EN_i, RegIMM_LATCH_EN => 
                           RegIMM_LATCH_EN_i, Reg_RD1_EN => en_RD1_i, RD1 => 
                           rd1_i, RD2 => rd2_i, B2_LATCH_EN => B2_EN_i, 
                           MUXA_SEL => MUXA_SEL_i, MUXB_SEL => MUXB_SEL_i, 
                           ALU_OUTREG_EN => ALU_OUTREG_EN_i, RETURN_REG_EN => 
                           RETURN_REG_EN_i, Reg_RD2_EN => en_RD2_i, DRAM_WE => 
                           net583, ALU_OUT2_SEL => sel_alu_ret_i, LMD_LATCH_EN 
                           => LMD_LATCH_EN_i, Alu_outreg2_en => 
                           Alu_outreg2_en_i, JUMP_en => JUMP_EN_i, PC_LATCH_EN 
                           => net584, Reg_RD3_EN => en_RD3_i, 
                           write_stop_if_branch => write_stop_if_branch_i, 
                           WB_MUX_SEL => WB_MUX_SEL_i, RF_WE => net585, 
                           WB_MUX_ADD_SEL => wb_mux_add_sel_i, WR => wr_cu);
   add_351 : DLX_IR_SIZE32_PC_SIZE32_DW01_add_0 port map( A(31) => npc2_31_port
                           , A(30) => npc2_30_port, A(29) => npc2_29_port, 
                           A(28) => npc2_28_port, A(27) => npc2_27_port, A(26) 
                           => npc2_26_port, A(25) => npc2_25_port, A(24) => 
                           npc2_24_port, A(23) => npc2_23_port, A(22) => 
                           npc2_22_port, A(21) => npc2_21_port, A(20) => 
                           npc2_20_port, A(19) => npc2_19_port, A(18) => 
                           npc2_18_port, A(17) => npc2_17_port, A(16) => 
                           npc2_16_port, A(15) => npc2_15_port, A(14) => 
                           npc2_14_port, A(13) => npc2_13_port, A(12) => 
                           npc2_12_port, A(11) => npc2_11_port, A(10) => 
                           npc2_10_port, A(9) => npc2_9_port, A(8) => 
                           npc2_8_port, A(7) => npc2_7_port, A(6) => 
                           npc2_6_port, A(5) => npc2_5_port, A(4) => 
                           npc2_4_port, A(3) => npc2_3_port, A(2) => 
                           npc2_2_port, A(1) => npc2_1_port, A(0) => 
                           npc2_0_port, B(31) => immediate_31_port, B(30) => 
                           immediate_30_port, B(29) => immediate_29_port, B(28)
                           => immediate_28_port, B(27) => immediate_27_port, 
                           B(26) => immediate_26_port, B(25) => 
                           immediate_25_port, B(24) => immediate_24_port, B(23)
                           => immediate_23_port, B(22) => immediate_22_port, 
                           B(21) => immediate_21_port, B(20) => 
                           immediate_20_port, B(19) => immediate_19_port, B(18)
                           => immediate_18_port, B(17) => immediate_17_port, 
                           B(16) => immediate_16_port, B(15) => 
                           immediate_15_port, B(14) => immediate_14_port, B(13)
                           => immediate_13_port, B(12) => immediate_12_port, 
                           B(11) => immediate_11_port, B(10) => 
                           immediate_10_port, B(9) => immediate_9_port, B(8) =>
                           immediate_8_port, B(7) => immediate_7_port, B(6) => 
                           immediate_6_port, B(5) => immediate_5_port, B(4) => 
                           immediate_4_port, B(3) => immediate_3_port, B(2) => 
                           immediate_2_port, B(1) => immediate_1_port, B(0) => 
                           immediate_0_port, CI => n1, SUM(31) => 
                           pc_jump_31_port, SUM(30) => pc_jump_30_port, SUM(29)
                           => pc_jump_29_port, SUM(28) => pc_jump_28_port, 
                           SUM(27) => pc_jump_27_port, SUM(26) => 
                           pc_jump_26_port, SUM(25) => pc_jump_25_port, SUM(24)
                           => pc_jump_24_port, SUM(23) => pc_jump_23_port, 
                           SUM(22) => pc_jump_22_port, SUM(21) => 
                           pc_jump_21_port, SUM(20) => pc_jump_20_port, SUM(19)
                           => pc_jump_19_port, SUM(18) => pc_jump_18_port, 
                           SUM(17) => pc_jump_17_port, SUM(16) => 
                           pc_jump_16_port, SUM(15) => pc_jump_15_port, SUM(14)
                           => pc_jump_14_port, SUM(13) => pc_jump_13_port, 
                           SUM(12) => pc_jump_12_port, SUM(11) => 
                           pc_jump_11_port, SUM(10) => pc_jump_10_port, SUM(9) 
                           => pc_jump_9_port, SUM(8) => pc_jump_8_port, SUM(7) 
                           => pc_jump_7_port, SUM(6) => pc_jump_6_port, SUM(5) 
                           => pc_jump_5_port, SUM(4) => pc_jump_4_port, SUM(3) 
                           => pc_jump_3_port, SUM(2) => pc_jump_2_port, SUM(1) 
                           => pc_jump_1_port, SUM(0) => pc_jump_0_port, CO => 
                           net43113);
   add_306 : DLX_IR_SIZE32_PC_SIZE32_DW01_add_1 port map( A(31) => PC_31_port, 
                           A(30) => PC_30_port, A(29) => PC_29_port, A(28) => 
                           PC_28_port, A(27) => PC_27_port, A(26) => PC_26_port
                           , A(25) => PC_25_port, A(24) => PC_24_port, A(23) =>
                           PC_23_port, A(22) => PC_22_port, A(21) => PC_21_port
                           , A(20) => PC_20_port, A(19) => PC_19_port, A(18) =>
                           PC_18_port, A(17) => PC_17_port, A(16) => PC_16_port
                           , A(15) => PC_15_port, A(14) => PC_14_port, A(13) =>
                           PC_13_port, A(12) => PC_12_port, A(11) => PC_11_port
                           , A(10) => PC_10_port, A(9) => PC_9_port, A(8) => 
                           PC_8_port, A(7) => PC_7_port, A(6) => PC_6_port, 
                           A(5) => PC_5_port, A(4) => PC_4_port, A(3) => 
                           PC_3_port, A(2) => PC_2_port, A(1) => PC_1_port, 
                           A(0) => PC_0_port, B(31) => n2, B(30) => n2, B(29) 
                           => n2, B(28) => n2, B(27) => n2, B(26) => n2, B(25) 
                           => n2, B(24) => n2, B(23) => n2, B(22) => n2, B(21) 
                           => n2, B(20) => n2, B(19) => n2, B(18) => n2, B(17) 
                           => n2, B(16) => n2, B(15) => n2, B(14) => n2, B(13) 
                           => n2, B(12) => n2, B(11) => n2, B(10) => n2, B(9) 
                           => n2, B(8) => n2, B(7) => n2, B(6) => n2, B(5) => 
                           n2, B(4) => n2, B(3) => n2, B(2) => X_Logic1_port, 
                           B(1) => X_Logic0_port, B(0) => X_Logic0_port, CI => 
                           n2, SUM(31) => in_NPC_31_port, SUM(30) => 
                           in_NPC_30_port, SUM(29) => in_NPC_29_port, SUM(28) 
                           => in_NPC_28_port, SUM(27) => in_NPC_27_port, 
                           SUM(26) => in_NPC_26_port, SUM(25) => in_NPC_25_port
                           , SUM(24) => in_NPC_24_port, SUM(23) => 
                           in_NPC_23_port, SUM(22) => in_NPC_22_port, SUM(21) 
                           => in_NPC_21_port, SUM(20) => in_NPC_20_port, 
                           SUM(19) => in_NPC_19_port, SUM(18) => in_NPC_18_port
                           , SUM(17) => in_NPC_17_port, SUM(16) => 
                           in_NPC_16_port, SUM(15) => in_NPC_15_port, SUM(14) 
                           => in_NPC_14_port, SUM(13) => in_NPC_13_port, 
                           SUM(12) => in_NPC_12_port, SUM(11) => in_NPC_11_port
                           , SUM(10) => in_NPC_10_port, SUM(9) => in_NPC_9_port
                           , SUM(8) => in_NPC_8_port, SUM(7) => in_NPC_7_port, 
                           SUM(6) => in_NPC_6_port, SUM(5) => in_NPC_5_port, 
                           SUM(4) => in_NPC_4_port, SUM(3) => in_NPC_3_port, 
                           SUM(2) => in_NPC_2_port, SUM(1) => in_NPC_1_port, 
                           SUM(0) => in_NPC_0_port, CO => net43112);
   U267 : AND2_X2 port map( A1 => Rst, A2 => n298, ZN => n168);
   U268 : INV_X2 port map( A => n298, ZN => jump_verified);
   U269 : NOR2_X1 port map( A1 => write_stop_if_branch_i, A2 => n297, ZN => 
                           wr_i);
   U270 : INV_X1 port map( A => wr_cu, ZN => n297);
   U271 : MUX2_X1 port map( A => npc2_0_port, B => out_NPC_0_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n296);
   U272 : MUX2_X1 port map( A => PC_31_port, B => PC_BUS_31_port, S => 
                           NPC1_LATCH_EN_i, Z => n295);
   U273 : MUX2_X1 port map( A => out_NPC_31_port, B => in_NPC_31_port, S => 
                           NPC1_LATCH_EN_i, Z => n294);
   U274 : MUX2_X1 port map( A => npc2_31_port, B => out_NPC_31_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n293);
   U275 : MUX2_X1 port map( A => out_NPC_0_port, B => in_NPC_0_port, S => 
                           NPC1_LATCH_EN_i, Z => n292);
   U276 : MUX2_X1 port map( A => out_NPC_1_port, B => in_NPC_1_port, S => 
                           NPC1_LATCH_EN_i, Z => n291);
   U277 : MUX2_X1 port map( A => npc2_1_port, B => out_NPC_1_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n290);
   U278 : MUX2_X1 port map( A => out_NPC_2_port, B => in_NPC_2_port, S => 
                           NPC1_LATCH_EN_i, Z => n289);
   U279 : MUX2_X1 port map( A => npc2_2_port, B => out_NPC_2_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n288);
   U280 : MUX2_X1 port map( A => out_NPC_3_port, B => in_NPC_3_port, S => 
                           NPC1_LATCH_EN_i, Z => n287);
   U281 : MUX2_X1 port map( A => npc2_3_port, B => out_NPC_3_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n286);
   U282 : MUX2_X1 port map( A => out_NPC_4_port, B => in_NPC_4_port, S => 
                           NPC1_LATCH_EN_i, Z => n285);
   U283 : MUX2_X1 port map( A => npc2_4_port, B => out_NPC_4_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n284);
   U284 : MUX2_X1 port map( A => out_NPC_5_port, B => in_NPC_5_port, S => 
                           NPC1_LATCH_EN_i, Z => n283);
   U285 : MUX2_X1 port map( A => npc2_5_port, B => out_NPC_5_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n282);
   U286 : MUX2_X1 port map( A => out_NPC_6_port, B => in_NPC_6_port, S => 
                           NPC1_LATCH_EN_i, Z => n281);
   U287 : MUX2_X1 port map( A => npc2_6_port, B => out_NPC_6_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n280);
   U288 : MUX2_X1 port map( A => out_NPC_7_port, B => in_NPC_7_port, S => 
                           NPC1_LATCH_EN_i, Z => n279);
   U289 : MUX2_X1 port map( A => npc2_7_port, B => out_NPC_7_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n278);
   U290 : MUX2_X1 port map( A => out_NPC_8_port, B => in_NPC_8_port, S => 
                           NPC1_LATCH_EN_i, Z => n277);
   U291 : MUX2_X1 port map( A => npc2_8_port, B => out_NPC_8_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n276);
   U292 : MUX2_X1 port map( A => out_NPC_9_port, B => in_NPC_9_port, S => 
                           NPC1_LATCH_EN_i, Z => n275);
   U293 : MUX2_X1 port map( A => npc2_9_port, B => out_NPC_9_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n274);
   U294 : MUX2_X1 port map( A => out_NPC_10_port, B => in_NPC_10_port, S => 
                           NPC1_LATCH_EN_i, Z => n273);
   U295 : MUX2_X1 port map( A => npc2_10_port, B => out_NPC_10_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n272);
   U296 : MUX2_X1 port map( A => out_NPC_11_port, B => in_NPC_11_port, S => 
                           NPC1_LATCH_EN_i, Z => n271);
   U297 : MUX2_X1 port map( A => npc2_11_port, B => out_NPC_11_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n270);
   U298 : MUX2_X1 port map( A => out_NPC_12_port, B => in_NPC_12_port, S => 
                           NPC1_LATCH_EN_i, Z => n269);
   U299 : MUX2_X1 port map( A => npc2_12_port, B => out_NPC_12_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n268);
   U300 : MUX2_X1 port map( A => out_NPC_13_port, B => in_NPC_13_port, S => 
                           NPC1_LATCH_EN_i, Z => n267);
   U301 : MUX2_X1 port map( A => npc2_13_port, B => out_NPC_13_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n266);
   U302 : MUX2_X1 port map( A => out_NPC_14_port, B => in_NPC_14_port, S => 
                           NPC1_LATCH_EN_i, Z => n265);
   U303 : MUX2_X1 port map( A => npc2_14_port, B => out_NPC_14_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n264);
   U304 : MUX2_X1 port map( A => out_NPC_15_port, B => in_NPC_15_port, S => 
                           NPC1_LATCH_EN_i, Z => n263);
   U305 : MUX2_X1 port map( A => npc2_15_port, B => out_NPC_15_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n262);
   U306 : MUX2_X1 port map( A => out_NPC_16_port, B => in_NPC_16_port, S => 
                           NPC1_LATCH_EN_i, Z => n261);
   U307 : MUX2_X1 port map( A => npc2_16_port, B => out_NPC_16_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n260);
   U308 : MUX2_X1 port map( A => out_NPC_17_port, B => in_NPC_17_port, S => 
                           NPC1_LATCH_EN_i, Z => n259);
   U309 : MUX2_X1 port map( A => npc2_17_port, B => out_NPC_17_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n258);
   U310 : MUX2_X1 port map( A => out_NPC_18_port, B => in_NPC_18_port, S => 
                           NPC1_LATCH_EN_i, Z => n257);
   U311 : MUX2_X1 port map( A => npc2_18_port, B => out_NPC_18_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n256);
   U312 : MUX2_X1 port map( A => out_NPC_19_port, B => in_NPC_19_port, S => 
                           NPC1_LATCH_EN_i, Z => n255);
   U313 : MUX2_X1 port map( A => npc2_19_port, B => out_NPC_19_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n254);
   U314 : MUX2_X1 port map( A => out_NPC_20_port, B => in_NPC_20_port, S => 
                           NPC1_LATCH_EN_i, Z => n253);
   U315 : MUX2_X1 port map( A => npc2_20_port, B => out_NPC_20_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n252);
   U316 : MUX2_X1 port map( A => out_NPC_21_port, B => in_NPC_21_port, S => 
                           NPC1_LATCH_EN_i, Z => n251);
   U317 : MUX2_X1 port map( A => npc2_21_port, B => out_NPC_21_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n250);
   U318 : MUX2_X1 port map( A => out_NPC_22_port, B => in_NPC_22_port, S => 
                           NPC1_LATCH_EN_i, Z => n249);
   U319 : MUX2_X1 port map( A => npc2_22_port, B => out_NPC_22_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n248);
   U320 : MUX2_X1 port map( A => out_NPC_23_port, B => in_NPC_23_port, S => 
                           NPC1_LATCH_EN_i, Z => n247);
   U321 : MUX2_X1 port map( A => npc2_23_port, B => out_NPC_23_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n246);
   U322 : MUX2_X1 port map( A => out_NPC_24_port, B => in_NPC_24_port, S => 
                           NPC1_LATCH_EN_i, Z => n245);
   U323 : MUX2_X1 port map( A => npc2_24_port, B => out_NPC_24_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n244);
   U324 : MUX2_X1 port map( A => out_NPC_25_port, B => in_NPC_25_port, S => 
                           NPC1_LATCH_EN_i, Z => n243);
   U325 : MUX2_X1 port map( A => npc2_25_port, B => out_NPC_25_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n242);
   U326 : MUX2_X1 port map( A => out_NPC_26_port, B => in_NPC_26_port, S => 
                           NPC1_LATCH_EN_i, Z => n241);
   U327 : MUX2_X1 port map( A => npc2_26_port, B => out_NPC_26_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n240);
   U328 : MUX2_X1 port map( A => out_NPC_27_port, B => in_NPC_27_port, S => 
                           NPC1_LATCH_EN_i, Z => n239);
   U329 : MUX2_X1 port map( A => npc2_27_port, B => out_NPC_27_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n238);
   U330 : MUX2_X1 port map( A => out_NPC_28_port, B => in_NPC_28_port, S => 
                           NPC1_LATCH_EN_i, Z => n237);
   U331 : MUX2_X1 port map( A => npc2_28_port, B => out_NPC_28_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n236);
   U332 : MUX2_X1 port map( A => out_NPC_29_port, B => in_NPC_29_port, S => 
                           NPC1_LATCH_EN_i, Z => n235);
   U333 : MUX2_X1 port map( A => npc2_29_port, B => out_NPC_29_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n234);
   U334 : MUX2_X1 port map( A => out_NPC_30_port, B => in_NPC_30_port, S => 
                           NPC1_LATCH_EN_i, Z => n233);
   U335 : MUX2_X1 port map( A => npc2_30_port, B => out_NPC_30_port, S => 
                           RegAluOpCodeGen_EN_i, Z => n232);
   U336 : MUX2_X1 port map( A => PC_0_port, B => PC_BUS_0_port, S => 
                           NPC1_LATCH_EN_i, Z => n231);
   U337 : MUX2_X1 port map( A => PC_1_port, B => PC_BUS_1_port, S => 
                           NPC1_LATCH_EN_i, Z => n230);
   U338 : MUX2_X1 port map( A => PC_2_port, B => PC_BUS_2_port, S => 
                           NPC1_LATCH_EN_i, Z => n229);
   U339 : MUX2_X1 port map( A => PC_3_port, B => PC_BUS_3_port, S => 
                           NPC1_LATCH_EN_i, Z => n228);
   U340 : MUX2_X1 port map( A => PC_4_port, B => PC_BUS_4_port, S => 
                           NPC1_LATCH_EN_i, Z => n227);
   U341 : MUX2_X1 port map( A => PC_5_port, B => PC_BUS_5_port, S => 
                           NPC1_LATCH_EN_i, Z => n226);
   U342 : MUX2_X1 port map( A => PC_6_port, B => PC_BUS_6_port, S => 
                           NPC1_LATCH_EN_i, Z => n225);
   U343 : MUX2_X1 port map( A => PC_7_port, B => PC_BUS_7_port, S => 
                           NPC1_LATCH_EN_i, Z => n224);
   U344 : MUX2_X1 port map( A => PC_8_port, B => PC_BUS_8_port, S => 
                           NPC1_LATCH_EN_i, Z => n223);
   U345 : MUX2_X1 port map( A => PC_9_port, B => PC_BUS_9_port, S => 
                           NPC1_LATCH_EN_i, Z => n222);
   U346 : MUX2_X1 port map( A => PC_10_port, B => PC_BUS_10_port, S => 
                           NPC1_LATCH_EN_i, Z => n221);
   U347 : MUX2_X1 port map( A => PC_11_port, B => PC_BUS_11_port, S => 
                           NPC1_LATCH_EN_i, Z => n220);
   U348 : MUX2_X1 port map( A => PC_12_port, B => PC_BUS_12_port, S => 
                           NPC1_LATCH_EN_i, Z => n219);
   U349 : MUX2_X1 port map( A => PC_13_port, B => PC_BUS_13_port, S => 
                           NPC1_LATCH_EN_i, Z => n218);
   U350 : MUX2_X1 port map( A => PC_14_port, B => PC_BUS_14_port, S => 
                           NPC1_LATCH_EN_i, Z => n217);
   U351 : MUX2_X1 port map( A => PC_15_port, B => PC_BUS_15_port, S => 
                           NPC1_LATCH_EN_i, Z => n216);
   U352 : MUX2_X1 port map( A => PC_16_port, B => PC_BUS_16_port, S => 
                           NPC1_LATCH_EN_i, Z => n215);
   U353 : MUX2_X1 port map( A => PC_17_port, B => PC_BUS_17_port, S => 
                           NPC1_LATCH_EN_i, Z => n214);
   U354 : MUX2_X1 port map( A => PC_18_port, B => PC_BUS_18_port, S => 
                           NPC1_LATCH_EN_i, Z => n213);
   U355 : MUX2_X1 port map( A => PC_19_port, B => PC_BUS_19_port, S => 
                           NPC1_LATCH_EN_i, Z => n212);
   U356 : MUX2_X1 port map( A => PC_20_port, B => PC_BUS_20_port, S => 
                           NPC1_LATCH_EN_i, Z => n211);
   U357 : MUX2_X1 port map( A => PC_21_port, B => PC_BUS_21_port, S => 
                           NPC1_LATCH_EN_i, Z => n210);
   U358 : MUX2_X1 port map( A => PC_22_port, B => PC_BUS_22_port, S => 
                           NPC1_LATCH_EN_i, Z => n209);
   U359 : MUX2_X1 port map( A => PC_23_port, B => PC_BUS_23_port, S => 
                           NPC1_LATCH_EN_i, Z => n208);
   U360 : MUX2_X1 port map( A => PC_24_port, B => PC_BUS_24_port, S => 
                           NPC1_LATCH_EN_i, Z => n207);
   U361 : MUX2_X1 port map( A => PC_25_port, B => PC_BUS_25_port, S => 
                           NPC1_LATCH_EN_i, Z => n206);
   U362 : MUX2_X1 port map( A => PC_26_port, B => PC_BUS_26_port, S => 
                           NPC1_LATCH_EN_i, Z => n205);
   U363 : MUX2_X1 port map( A => PC_27_port, B => PC_BUS_27_port, S => 
                           NPC1_LATCH_EN_i, Z => n204);
   U364 : MUX2_X1 port map( A => PC_28_port, B => PC_BUS_28_port, S => 
                           NPC1_LATCH_EN_i, Z => n203);
   U365 : MUX2_X1 port map( A => PC_29_port, B => PC_BUS_29_port, S => 
                           NPC1_LATCH_EN_i, Z => n202);
   U366 : MUX2_X1 port map( A => PC_30_port, B => PC_BUS_30_port, S => 
                           NPC1_LATCH_EN_i, Z => n201);
   U367 : MUX2_X1 port map( A => IR_7_port, B => iram_Dout(7), S => 
                           NPC1_LATCH_EN_i, Z => n200);
   U368 : MUX2_X1 port map( A => IR_5_port, B => iram_Dout(5), S => 
                           NPC1_LATCH_EN_i, Z => n199);
   U369 : MUX2_X1 port map( A => IR_3_port, B => iram_Dout(3), S => 
                           NPC1_LATCH_EN_i, Z => n198);
   U370 : MUX2_X1 port map( A => IR_31_port, B => iram_Dout(31), S => 
                           NPC1_LATCH_EN_i, Z => n197);
   U371 : MUX2_X1 port map( A => IR_29_port, B => iram_Dout(29), S => 
                           NPC1_LATCH_EN_i, Z => n196);
   U372 : MUX2_X1 port map( A => IR_1_port, B => iram_Dout(1), S => 
                           NPC1_LATCH_EN_i, Z => n195);
   U373 : MUX2_X1 port map( A => IR_26_port, B => iram_Dout(26), S => 
                           NPC1_LATCH_EN_i, Z => n194);
   U374 : MUX2_X1 port map( A => IR_24_port, B => iram_Dout(24), S => 
                           NPC1_LATCH_EN_i, Z => n193);
   U375 : MUX2_X1 port map( A => IR_22_port, B => iram_Dout(22), S => 
                           NPC1_LATCH_EN_i, Z => n192);
   U376 : MUX2_X1 port map( A => IR_20_port, B => iram_Dout(20), S => 
                           NPC1_LATCH_EN_i, Z => n191);
   U377 : MUX2_X1 port map( A => IR_18_port, B => iram_Dout(18), S => 
                           NPC1_LATCH_EN_i, Z => n190);
   U378 : MUX2_X1 port map( A => IR_17_port, B => iram_Dout(17), S => 
                           NPC1_LATCH_EN_i, Z => n189);
   U379 : MUX2_X1 port map( A => IR_15_port, B => iram_Dout(15), S => 
                           NPC1_LATCH_EN_i, Z => n188);
   U380 : MUX2_X1 port map( A => IR_13_port, B => iram_Dout(13), S => 
                           NPC1_LATCH_EN_i, Z => n187);
   U381 : MUX2_X1 port map( A => IR_11_port, B => iram_Dout(11), S => 
                           NPC1_LATCH_EN_i, Z => n186);
   U382 : MUX2_X1 port map( A => IR_9_port, B => iram_Dout(9), S => 
                           NPC1_LATCH_EN_i, Z => n185);
   U383 : MUX2_X1 port map( A => IR_8_port, B => iram_Dout(8), S => 
                           NPC1_LATCH_EN_i, Z => n184);
   U384 : MUX2_X1 port map( A => IR_10_port, B => iram_Dout(10), S => 
                           NPC1_LATCH_EN_i, Z => n183);
   U385 : MUX2_X1 port map( A => IR_12_port, B => iram_Dout(12), S => 
                           NPC1_LATCH_EN_i, Z => n182);
   U386 : MUX2_X1 port map( A => IR_14_port, B => iram_Dout(14), S => 
                           NPC1_LATCH_EN_i, Z => n181);
   U387 : MUX2_X1 port map( A => IR_16_port, B => iram_Dout(16), S => 
                           NPC1_LATCH_EN_i, Z => n180);
   U388 : MUX2_X1 port map( A => IR_0_port, B => iram_Dout(0), S => 
                           NPC1_LATCH_EN_i, Z => n179);
   U389 : MUX2_X1 port map( A => IR_19_port, B => iram_Dout(19), S => 
                           NPC1_LATCH_EN_i, Z => n178);
   U390 : MUX2_X1 port map( A => IR_21_port, B => iram_Dout(21), S => 
                           NPC1_LATCH_EN_i, Z => n177);
   U391 : MUX2_X1 port map( A => IR_23_port, B => iram_Dout(23), S => 
                           NPC1_LATCH_EN_i, Z => n176);
   U392 : MUX2_X1 port map( A => IR_25_port, B => iram_Dout(25), S => 
                           NPC1_LATCH_EN_i, Z => n175);
   U393 : MUX2_X1 port map( A => IR_27_port, B => iram_Dout(27), S => 
                           NPC1_LATCH_EN_i, Z => n174);
   U394 : MUX2_X1 port map( A => IR_28_port, B => iram_Dout(28), S => 
                           NPC1_LATCH_EN_i, Z => n173);
   U395 : MUX2_X1 port map( A => IR_30_port, B => iram_Dout(30), S => 
                           NPC1_LATCH_EN_i, Z => n172);
   U396 : MUX2_X1 port map( A => IR_2_port, B => iram_Dout(2), S => 
                           NPC1_LATCH_EN_i, Z => n171);
   U397 : MUX2_X1 port map( A => IR_4_port, B => iram_Dout(4), S => 
                           NPC1_LATCH_EN_i, Z => n170);
   U398 : MUX2_X1 port map( A => IR_6_port, B => iram_Dout(6), S => 
                           NPC1_LATCH_EN_i, Z => n169);
   U399 : NOR2_X1 port map( A1 => JUMP_EN_i, A2 => comp_branch_dp, ZN => n298);

end SYN_dlx_rtl;
