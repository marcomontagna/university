LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
ENTITY MUX_10_to_1 IS
PORT(
SEL	: IN STD_LOGIC_VECTOR(3 DOWNTO 0);	--segnale di enable, reset e clock
DATA_0, DATA_1, DATA_2,DATA_3,DATA_4,DATA_5	:	IN STD_LOGIC;	--dato in ingresso
DATA_6, DATA_7, DATA_8, DATA_9 :	IN STD_LOGIC;	--dato in ingresso
DATA_OUT	:	OUT STD_LOGIC --dato in uscita
);
END ENTITY MUX_10_to_1;
ARCHITECTURE BEHAVIOR OF MUX_10_to_1 IS
BEGIN
WITH SEL SELECT DATA_OUT<=
DATA_0 WHEN "0000",
DATA_1 WHEN "0001",
DATA_2 WHEN "0010",
DATA_3 WHEN "0011",
DATA_4 WHEN "0100",
DATA_5 WHEN "0101",
DATA_6 WHEN "0110",
DATA_7 WHEN "0111",
DATA_8 WHEN "1000",
DATA_9 WHEN "1001",
DATA_0 WHEN OTHERS;
END BEHAVIOR;