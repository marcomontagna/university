library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned.all;
use IEEE.std_logic_arith.all;
use work.globals.all;

entity ALU is
  generic (N : integer := NumBit);
  port 	 ( AluOpCode: IN std_logic_vector(2 downto 0); -- selctor of which output operation choose (add/sub or and/or/xor or srl/sll)
	   CompareOpCode: in std_logic_vector(3 downto 0); --selection of type of compare operation CompareOpCode(3)->beqz
--												    CompareOpCode(2)->bnez
-- 												    CompareOpCode(1)->sge
--												    CompareOpCode(0)->sne   
	   Add_subn: in std_logic; --id add=0 if sub =1
	   ShiftOpCode:in std_logic_vector(2 downto 0);--specify the type of op for the shifter component: ShiftOpCode(2)->logic_arith
--     													ShiftOpCode(1)->LEFT_RIGHT
--													ShiftOpCode(0)->shift_rotate
								
           DATA1, DATA2: IN std_logic_vector(N-1 downto 0);
           OUTALU: OUT std_logic_vector(N-1 downto 0);
           return_address: buffer std_logic_vector(N-1 downto 0);
	   CompBranch: out std_logic);
end ALU;

architecture BEHAVIOR of ALU is

component SHIFTER_GENERIC is
	generic(N: integer);
	port(	A: in std_logic_vector(N-1 downto 0);
		B: in std_logic_vector(4 downto 0);
		LOGIC_ARITH: in std_logic;	-- 1 = logic, 0 = arith
		LEFT_RIGHT: in std_logic;	-- 1 = left, 0 = right
		SHIFT_ROTATE: in std_logic;	-- 1 = shift, 0 = rotate
		OUTPUT: out std_logic_vector(N-1 downto 0)
	);
end component;

component operatore_logic is 
    generic (REG_SIZE: INTEGER :=32);
	Port(	
			A:	In	std_logic_vector(REG_SIZE-1 downto 0);
			B:	In	std_logic_vector(REG_SIZE-1 downto 0);
			OUT_LOGIC_AND:	Out	std_logic_vector(REG_SIZE-1 downto 0);
			OUT_LOGIC_OR:	Out	std_logic_vector(REG_SIZE-1 downto 0);
			OUT_LOGIC_XOR:	Out	std_logic_vector(REG_SIZE-1 downto 0)
		   );
end component; 


component p4_adder is
  generic (
         N : integer :=32 ;
	 N_carry : integer :=4 );
	 
	 port( A: in std_logic_vector( N-1 downto 0);
		B :in std_logic_vector( N-1 downto 0);
		Cin : in std_logic;
		SUM : out std_logic_vector(N-1 downto 0));
end component;

component compare is
generic (N: integer:=32);
port(    num1 : in std_logic_vector(N-1 downto 0);  --input 1
         num2 : in std_logic_vector(N-1 downto 0);  --input 2
         less : out std_logic;   -- indicates first number is small
         equal: out std_logic;   -- both are equal
         greater:out std_logic    -- indicates first number is bigger
);
end component;

component MUX_6to1  
	generic (n: integer:=32);
	Port (	
		A:	In	std_logic_vector(n-1 downto 0); 
		B:	In	std_logic_vector(n-1 downto 0);
		C:	In	std_logic_vector(n-1 downto 0);
		D:	In	std_logic_vector(n-1 downto 0); 
		E:	In	std_logic_vector(n-1 downto 0);
		F:	In	std_logic_vector(n-1 downto 0);
		S:	In	std_logic_vector(2 downto 0);
		Y:	Out	std_logic_vector(n-1 downto 0));
end component;


component MUX_2to1 is 
	generic (n: integer:=32);
	Port (	
		A:	In	std_logic_vector(n-1 downto 0); 
		B:	In	std_logic_vector(n-1 downto 0);
		S:	In	std_logic;
		Y:	Out	std_logic_vector(n-1 downto 0));
end component ;

component RCA_GEN is
  generic (
    NBIT  : INTEGER := 16);
  port (
    A  : in     std_logic_vector(NBIT-1 downto 0);
    B  : in     std_logic_vector(NBIT -1 downto 0);
    Ci : in     std_logic;
    S  : buffer std_logic_vector(NBIT-1 downto 0);
    Co : out    std_logic);
end component;


signal AND_OUT, OR_OUT, XOR_OUT, comp_out, one_32bits, zero_32bits, four_32bits: std_logic_vector(NumBit-1 downto 0);

signal shift_out, add_sub_out: std_logic_vector(NUmBIt-1 downto 0);

signal comp_less, comp_eq, comp_greater, sge_verified, sne_verified, beqz_verified, bnez_verified, sel_mux_comp_out: std_logic;

begin

four_32bits(31 downto 3)<=(others=>'0');
four_32bits(2 downto 0)<="100";

adder4 : RCA_GEN generic map (32) --registro per return address (operazione jal)
port map(DATA1, four_32bits, '0', return_address, open); --prima c'�era data2

shifter: SHIFTER_GENERIC generic map(NumBit)
port map(DATA1, DATA2(4 downto 0), ShiftOpCode(2),  ShiftOpCode(1),  ShiftOpCode(0), shift_out); --31 27

logic_operations: operatore_logic generic map(N)
port map(DATA1, DATA2, AND_OUT, OR_OUT, XOR_OUT);

adder_sub: p4_adder generic map (32, 4)
port map(DATA1, DATA2, add_subn, add_sub_out);

comp: compare generic map (32)
port map(DATA1, DATA2, COMP_LESS, COMP_EQ, COMP_GREATER);

sge_verified<=(COMP_EQ OR COMP_GREATER) AND CompareOpCode(1);
sne_verified<=(NOT(COMP_EQ) AND CompareOpCode(0));
sel_mux_comp_out<= sne_verified or sge_verified;

one_32bits(31 downto 1)<=(others=>'0');
one_32bits(0)<='1';
zero_32bits<=(others=>'0');

mux_comp: mux_2to1 generic map (32)
port map(zero_32bits, one_32bits, sel_mux_comp_out, comp_out);

beqz_verified<=CompareOpCode(3) and COMP_EQ;
bnez_verified<=CompareOpCode(2) and NOT(COMP_EQ);

CompBranch<= bnez_verified or beqz_verified;

mux_alu_out: MUX_6to1 generic map (32)
port map (add_sub_out, and_out, or_out, xor_out, comp_out, shift_out, AluOpCode, outALU);
 
end BEHAVIOR;
